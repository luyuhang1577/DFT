1    20    0    1    0
1    311    0    1    0
1    45    0    1    0
1    107    0    1    0
1    41    0    1    0
1    179    0    1    0
1    116    0    1    0
1    97    0    1    0
1    77    0    1    0
1    132    0    1    0
1    169    0    1    0
1    274    0    1    0
1    33    0    1    0
1    68    0    1    0
1    244    0    1    0
1    213    0    1    0
1    283    0    1    0
1    190    0    1    0
1    250    0    1    0
1    124    0    1    0
1    329    0    1    0
1    87    0    1    0
1    128    0    1    0
1    222    0    1    0
1    232    0    1    0
1    226    0    1    0
1    13    0    1    0
1    264    0    1    0
1    200    0    1    0
1    150    0    1    0
1    159    0    1    0
1    326    0    1    0
1    317    0    1    0
1    125    0    1    0
1    238    0    1    0
1    322    0    1    0
1    294    0    1    0
1    137    0    1    0
1    1    0    1    0
1    1698    0    1    0
1    257    0    1    0
1    143    0    1    0
1    50    0    1    0
1    343    0    1    0
1    270    0    1    0
1    330    0    1    0
1    2897    0    1    0
1    223    0    1    0
1    303    0    1    0
1    58    0    1    0
2    432    1    50
0    442    5    1    1    50
2    447    1    58
0    456    5    1    1    58
2    460    1    68
0    463    5    1    1    68
2    467    1    68
2    476    1    77
0    479    5    1    1    77
2    483    1    77
2    492    1    87
0    501    5    1    1    87
2    504    1    97
0    513    5    1    1    97
2    517    1    107
0    526    5    1    1    107
2    530    1    116
0    540    5    1    1    116
0    587    3    1    2    257    264
0    704    5    1    1    1
2    707    1    1
0    714    5    1    1    1
2    717    1    13
0    724    5    1    1    13
0    731    7    1    2    13    20
0    732    5    1    1    20
2    736    1    20
0    741    5    1    1    20
0    758    5    1    1    33
2    776    1    33
0    780    5    1    1    33
0    788    7    1    2    33    41
0    791    5    1    1    41
0    798    3    1    2    41    45
2    799    1    45
0    802    5    1    1    45
0    826    5    1    1    50
2    828    1    58
0    831    5    1    1    58
2    833    1    68
0    836    5    1    1    68
2    839    1    87
0    842    5    1    1    87
2    845    1    97
0    848    5    1    1    97
0    851    5    1    1    107
2    890    1    1
2    898    1    68
2    907    1    107
0    1032    5    1    1    20
2    1035    1    190
0    1048    5    1    1    200
0    1049    7    1    2    20    200
0    1050    6    1    2    20    200
0    1051    7    1    2    20    179
0    1540    5    1    1    20
0    1699    3    1    2    1698    33
0    1826    6    1    2    1    13
0    1827    6    1    3    1    20    33
0    1828    5    1    1    20
0    2051    5    1    1    33
2    2478    1    179
0    2865    5    1    1    213
2    2868    1    343
2    2931    1    226
2    2934    1    232
2    2939    1    238
2    2942    1    244
2    2947    1    250
2    2950    1    257
2    2957    1    264
2    2960    1    270
2    3007    1    50
2    3079    1    58
2    3087    1    58
2    3095    1    97
2    3103    1    97
2    3419    1    330
0    588    7    1    2    250    587
0    759    3    1    2    758    20
0    1541    3    1    2    1540    169
0    1772    5    1    1    731
0    1829    3    1    2    1828    1
0    1834    7    1    2    1826    1827
0    2052    3    1    2    2051    1
0    625    7    1    3    826    831    836
0    545    6    1    2    226    432
0    546    6    1    2    232    447
0    547    6    1    2    238    467
0    548    6    1    2    244    483
0    549    6    1    2    250    492
0    550    6    1    2    257    504
0    551    6    1    2    264    517
0    552    6    1    2    270    530
0    2937    5    1    1    2931
0    2938    5    1    1    2934
0    2945    5    1    1    2939
0    2946    5    1    1    2942
0    621    6    1    2    456    463
0    626    6    1    2    513    526
0    635    6    1    2    460    476
2    636    1    442
0    3085    5    1    1    3079
0    3101    5    1    1    3095
2    657    1    802
2    675    1    802
2    721    1    717
2    784    1    780
2    794    1    791
0    807    7    1    2    714    798
0    816    7    1    3    714    799    791
0    823    7    1    2    704    799
0    860    7    1    3    707    724    736
0    861    6    1    3    707    724    736
0    864    6    1    2    707    724
2    893    1    890
0    896    6    1    3    717    732    45
0    897    6    1    3    826    831    836
0    3093    5    1    1    3087
0    905    7    1    3    842    848    851
0    906    6    1    3    842    848    851
0    3109    5    1    1    3103
0    973    5    1    1    741
0    980    5    1    1    741
0    987    5    1    1    741
0    994    5    1    1    741
0    1001    5    1    1    741
0    1008    5    1    1    741
0    1015    5    1    1    741
0    1022    5    1    1    741
0    1038    3    1    2    1032    1035
0    1043    4    1    2    1032    1035
2    1054    1    1051
0    1057    5    1    1    1051
2    1512    1    776
2    1681    1    780
0    1717    5    1    1    1699
0    1724    5    1    1    1699
0    1731    5    1    1    1699
0    1738    5    1    1    1699
0    1745    5    1    1    1699
0    1752    5    1    1    1699
0    1759    5    1    1    1699
0    1766    5    1    1    1699
0    1773    3    1    2    1    1772
0    1790    5    1    1    788
0    1808    5    1    1    788
0    2278    7    1    3    704    717    732
0    2481    5    1    1    2478
0    3425    5    1    1    3419
0    2871    3    1    2    2865    2868
0    2874    4    1    2    2865    2868
0    2953    5    1    1    2947
0    2954    5    1    1    2950
0    2963    5    1    1    2957
0    2964    5    1    1    2960
2    3010    1    456
0    3013    5    1    1    3007
2    3017    1    463
2    3020    1    479
2    3027    1    501
2    3030    1    513
2    3037    1    526
2    3040    1    540
2    3082    1    898
2    3090    1    898
2    3098    1    907
2    3106    1    907
0    352    6    1    2    479    625
0    553    7    1    4    545    546    547    548
0    554    7    1    4    549    550    551    552
0    555    6    1    2    2934    2937
0    556    6    1    2    2931    2938
0    560    6    1    2    2942    2945
0    561    6    1    2    2939    2946
0    650    7    1    2    432    621
0    956    7    1    2    890    896
0    974    5    1    1    759
0    975    7    1    2    741    759
0    976    7    1    2    897    973
0    981    5    1    1    759
0    982    7    1    2    741    759
0    988    5    1    1    759
0    989    7    1    2    741    759
0    990    7    1    2    836    987
0    995    5    1    1    759
0    996    7    1    2    741    759
0    997    7    1    2    77    994
0    1002    5    1    1    759
0    1003    7    1    2    741    759
0    1004    7    1    2    906    1001
0    1009    5    1    1    759
0    1010    7    1    2    741    759
0    1016    5    1    1    759
0    1017    7    1    2    741    759
0    1018    7    1    2    851    1015
0    1023    5    1    1    759
0    1024    7    1    2    741    759
0    1025    7    1    2    116    1022
0    1720    7    1    2    222    1717
0    1727    7    1    2    223    1724
0    1734    7    1    2    226    1731
0    1741    7    1    2    232    1738
0    1748    7    1    2    238    1745
0    1755    7    1    2    244    1752
0    1762    7    1    2    250    1759
0    1769    7    1    2    257    1766
0    1791    7    1    3    1    13    1790
0    1809    7    1    3    1    13    1808
0    1851    5    1    1    1834
0    1901    5    1    1    1834
0    1952    5    1    1    1834
0    2002    5    1    1    1834
0    2057    5    1    1    1834
0    2109    5    1    1    1834
0    2162    5    1    1    1834
0    2214    5    1    1    1834
0    2955    6    1    2    2950    2953
0    2956    6    1    2    2947    2954
0    2965    6    1    2    2960    2963
0    2966    6    1    2    2957    2964
3    353    5    1    1    352
0    354    7    1    2    87    626
0    557    6    1    2    555    556
0    562    6    1    2    560    561
0    586    6    1    2    553    554
0    630    7    1    2    540    905
0    634    6    1    2    540    905
0    639    5    1    1    636
0    642    6    1    2    3082    3085
0    3086    5    1    1    3082
0    644    7    1    2    460    636
0    646    6    1    2    3098    3101
0    3102    5    1    1    3098
0    654    6    1    2    87    626
0    660    5    1    1    657
0    678    5    1    1    675
0    804    6    1    2    860    776
0    806    6    1    2    860    780
0    855    6    1    3    707    721    736
0    867    6    1    4    707    724    736    794
0    903    6    1    2    3090    3093
0    3094    5    1    1    3090
0    912    6    1    2    3106    3109
0    3110    5    1    1    3106
0    915    5    1    1    861
0    927    5    1    1    893
0    941    5    1    1    864
0    977    7    1    2    828    974
0    978    7    1    2    150    975
0    984    7    1    2    833    981
0    985    7    1    2    159    982
0    991    7    1    2    77    988
0    992    7    1    2    50    989
0    998    7    1    2    839    995
0    999    7    1    2    828    996
0    1005    7    1    2    845    1002
0    1006    7    1    2    833    1003
0    1012    7    1    2    107    1009
0    1013    7    1    2    77    1010
0    1019    7    1    2    116    1016
0    1020    7    1    2    839    1017
0    1026    7    1    2    283    1023
0    1027    7    1    2    845    1024
0    1060    7    1    2    200    1054
0    1063    7    1    2    1048    1054
0    1066    7    1    2    1049    1057
0    1069    7    1    2    1050    1057
0    1527    6    1    2    784    794
0    1530    6    1    2    776    794
0    1542    6    1    3    707    721    1541
0    1563    6    1    3    724    732    784
0    1572    6    1    2    724    784
0    1581    5    1    1    1512
0    1585    5    1    1    1512
0    1589    5    1    1    1512
0    1593    5    1    1    1512
0    1597    5    1    1    1512
0    1601    5    1    1    1512
0    1605    5    1    1    1512
0    1716    5    1    1    1681
0    1718    7    1    2    1681    1699
0    1723    5    1    1    1681
0    1725    7    1    2    1681    1699
0    1730    5    1    1    1681
0    1732    7    1    2    1681    1699
0    1737    5    1    1    1681
0    1739    7    1    2    1681    1699
0    1744    5    1    1    1681
0    1746    7    1    2    1681    1699
0    1751    5    1    1    1681
0    1753    7    1    2    1681    1699
0    1758    5    1    1    1681
0    1760    7    1    2    1681    1699
0    1765    5    1    1    1681
0    1767    7    1    2    1681    1699
0    1852    7    1    2    1834    1773
0    1856    4    1    2    50    1773
0    1870    5    1    1    807
0    1902    7    1    2    1834    1773
0    1906    4    1    2    58    1773
0    1920    5    1    1    807
0    1953    7    1    2    1834    1773
0    1957    4    1    2    68    1773
0    1971    5    1    1    807
0    2003    7    1    2    1834    1773
0    2007    4    1    2    77    1773
0    2021    5    1    1    807
0    2058    7    1    2    1834    1773
0    2062    4    1    2    87    1773
0    2076    5    1    1    823
0    2110    7    1    2    1834    1773
0    2114    4    1    2    97    1773
0    2128    5    1    1    816
0    2163    7    1    2    1834    1773
0    2167    4    1    2    107    1773
0    2181    5    1    1    816
0    2215    7    1    2    1834    1773
0    2219    4    1    2    116    1773
0    2233    5    1    1    816
0    2285    7    1    2    2278    213
0    2288    6    1    2    2278    213
0    2289    7    1    3    2278    213    343
0    2293    6    1    3    2278    213    343
0    2298    7    1    3    2278    213    343
0    2302    6    1    3    2278    213    343
2    2877    1    2874
0    2983    6    1    2    2955    2956
0    2986    6    1    2    2965    2966
0    3014    5    1    1    3010
0    3015    6    1    2    3010    3013
0    3023    5    1    1    3017
0    3024    5    1    1    3020
0    3033    5    1    1    3027
0    3034    5    1    1    3030
0    3043    5    1    1    3037
0    3044    5    1    1    3040
3    355    5    1    1    354
0    643    6    1    2    3079    3086
0    647    6    1    2    3095    3102
0    680    7    1    2    650    675
0    904    6    1    2    3087    3094
0    913    6    1    2    3103    3110
0    920    7    1    2    588    915
0    979    3    1    3    976    977    978
0    993    3    1    3    990    991    992
0    1000    3    1    3    997    998    999
0    1007    3    1    3    1004    1005    1006
0    1021    3    1    3    1018    1019    1020
0    1028    3    1    3    1025    1026    1027
0    1719    7    1    2    77    1716
0    1721    7    1    2    223    1718
0    1726    7    1    2    87    1723
0    1728    7    1    2    226    1725
0    1733    7    1    2    97    1730
0    1735    7    1    2    232    1732
0    1740    7    1    2    107    1737
0    1742    7    1    2    238    1739
0    1747    7    1    2    116    1744
0    1749    7    1    2    244    1746
0    1754    7    1    2    283    1751
0    1756    7    1    2    250    1753
0    1761    7    1    2    294    1758
0    1763    7    1    2    257    1760
0    1768    7    1    2    303    1765
0    1770    7    1    2    264    1767
2    1794    1    1791
0    1799    5    1    1    1791
2    1812    1    1809
0    1817    5    1    1    1809
0    1859    7    1    3    50    1829    1852
0    1909    7    1    3    58    1829    1902
0    1960    7    1    3    68    1829    1953
0    2010    7    1    3    77    1829    2003
0    2065    7    1    3    87    2052    2058
0    2117    7    1    3    97    2052    2110
0    2170    7    1    3    107    2052    2163
0    2222    7    1    3    116    2052    2215
0    2678    5    1    1    956
0    2697    5    1    1    956
0    2716    5    1    1    956
0    2733    5    1    1    956
0    2751    5    1    1    956
0    2768    5    1    1    956
0    2785    5    1    1    956
0    2802    5    1    1    956
0    3016    6    1    2    3007    3014
0    3025    6    1    2    3020    3023
0    3026    6    1    2    3017    3024
0    3035    6    1    2    3030    3033
0    3036    6    1    2    3027    3034
0    3045    6    1    2    3040    3043
0    3046    6    1    2    3037    3044
0    2989    5    1    1    2983
0    2990    5    1    1    2986
0    610    5    1    1    804
0    613    7    1    2    804    806
0    616    5    1    1    806
0    640    6    1    2    642    643
0    648    6    1    2    646    647
0    655    7    1    4    630    635    442    58
0    665    5    1    1    804
0    668    7    1    2    804    806
0    671    5    1    1    806
0    683    5    1    1    804
0    685    5    1    1    806
0    688    7    1    2    804    806
0    694    5    1    1    804
0    696    5    1    1    806
0    699    7    1    2    804    806
2    870    1    867
2    887    1    867
0    901    6    1    2    903    904
0    910    6    1    2    912    913
0    914    5    1    1    855
0    916    7    1    2    855    861
0    942    5    1    1    855
0    943    7    1    2    864    855
0    1072    6    1    2    1043    1069
0    1084    6    1    2    1043    1066
0    1096    6    1    2    1038    1069
0    1108    6    1    2    1038    1066
0    1120    6    1    2    1043    1063
0    1132    6    1    2    1043    1060
0    1144    6    1    2    1038    1063
0    1156    6    1    2    1038    1060
0    1533    5    1    1    1527
0    1534    5    1    1    1530
0    1535    7    1    2    1527    1530
2    1545    1    1542
2    1554    1    1542
0    1610    5    1    1    1572
0    1619    5    1    1    1572
0    1628    5    1    1    1572
0    1637    5    1    1    1572
0    1646    5    1    1    1563
0    1655    5    1    1    1563
0    1664    5    1    1    1563
0    1673    5    1    1    1563
0    1722    3    1    3    1719    1720    1721
0    1729    3    1    3    1726    1727    1728
0    1736    3    1    3    1733    1734    1735
0    1743    3    1    3    1740    1741    1742
0    1750    3    1    3    1747    1748    1749
0    1757    3    1    3    1754    1755    1756
0    1764    3    1    3    1761    1762    1763
0    1771    3    1    3    1768    1769    1770
0    1853    7    1    2    979    1851
0    1954    7    1    2    993    1952
0    2004    7    1    2    1000    2002
0    2059    7    1    2    1007    2057
0    2164    7    1    2    1021    2162
0    2216    7    1    2    1028    2214
2    2485    1    2293
0    2900    7    1    2    2877    2897
0    2903    6    1    2    2877    2897
2    2967    1    557
2    2970    1    562
2    2975    1    557
2    2978    1    562
0    3047    6    1    2    3015    3016
0    3050    6    1    2    3025    3026
0    3055    6    1    2    3035    3036
0    3058    6    1    2    3045    3046
0    574    6    1    2    2986    2989
0    575    6    1    2    2983    2990
0    617    7    1    2    501    613
0    641    7    1    3    640    476    639
0    649    7    1    2    530    648
0    662    7    1    2    655    657
0    672    7    1    2    513    668
0    690    7    1    2    654    685
0    691    7    1    2    540    688
0    701    7    1    2    634    696
0    702    7    1    2    526    699
0    902    5    1    1    901
0    911    5    1    1    910
0    917    7    1    2    650    914
0    923    7    1    2    586    916
0    1538    7    1    2    442    1535
0    1871    7    1    3    1817    226    1870
0    1872    7    1    3    1817    274    807
0    1873    7    1    2    1812    1722
0    1921    7    1    3    1817    232    1920
0    1922    7    1    3    1817    274    807
0    1923    7    1    2    1812    1729
0    1972    7    1    3    1817    238    1971
0    1973    7    1    3    1817    274    807
0    1974    7    1    2    1812    1736
0    2022    7    1    3    1817    244    2021
0    2023    7    1    3    1817    274    807
0    2024    7    1    2    1812    1743
0    2077    7    1    3    1799    250    2076
0    2078    7    1    3    1799    274    823
0    2079    7    1    2    1794    1750
0    2129    7    1    3    1799    257    2128
0    2130    7    1    3    1799    274    816
0    2131    7    1    2    1794    1757
0    2182    7    1    3    1799    264    2181
0    2183    7    1    3    1799    274    816
0    2184    7    1    2    1794    1764
0    2234    7    1    3    1799    270    2233
0    2235    7    1    3    1799    274    816
0    2236    7    1    2    1794    1771
0    2973    5    1    1    2967
0    2974    5    1    1    2970
0    2981    5    1    1    2975
0    2982    5    1    1    2978
0    576    6    1    2    574    575
0    3053    5    1    1    3047
0    3054    5    1    1    3050
0    3061    5    1    1    3055
0    3062    5    1    1    3058
0    645    3    1    2    641    644
0    926    5    1    1    887
0    928    7    1    2    887    893
0    947    7    1    2    649    942
0    983    7    1    2    902    980
0    1011    7    1    2    911    1008
2    1075    1    1072
2    1087    1    1084
2    1099    1    1096
2    1111    1    1108
2    1123    1    1120
2    1135    1    1132
2    1147    1    1144
2    1159    1    1156
2    1168    1    1072
2    1177    1    1084
2    1186    1    1096
2    1195    1    1108
2    1204    1    1120
2    1213    1    1132
2    1222    1    1144
2    1231    1    1156
0    1609    5    1    1    1545
0    1611    7    1    2    1545    1572
0    1618    5    1    1    1545
0    1620    7    1    2    1545    1572
0    1627    5    1    1    1545
0    1629    7    1    2    1545    1572
0    1636    5    1    1    1545
0    1638    7    1    2    1545    1572
0    1645    5    1    1    1554
0    1647    7    1    2    1554    1563
0    1654    5    1    1    1554
0    1656    7    1    2    1554    1563
0    1663    5    1    1    1554
0    1665    7    1    2    1554    1563
0    1672    5    1    1    1554
0    1674    7    1    2    1554    1563
0    1862    3    1    3    1853    1856    1859
0    1866    4    1    3    1853    1856    1859
0    1874    3    1    3    1871    1872    1873
0    1924    3    1    3    1921    1922    1923
0    1963    3    1    3    1954    1957    1960
0    1967    4    1    3    1954    1957    1960
0    1975    3    1    3    1972    1973    1974
0    2013    3    1    3    2004    2007    2010
0    2017    4    1    3    2004    2007    2010
0    2025    3    1    3    2022    2023    2024
0    2068    3    1    3    2059    2062    2065
0    2072    4    1    3    2059    2062    2065
0    2080    3    1    3    2077    2078    2079
0    2132    3    1    3    2129    2130    2131
0    2173    3    1    3    2164    2167    2170
0    2177    4    1    3    2164    2167    2170
0    2185    3    1    3    2182    2183    2184
0    2225    3    1    3    2216    2219    2222
0    2229    4    1    3    2216    2219    2222
0    2237    3    1    3    2234    2235    2236
0    2488    5    1    1    2485
0    2679    5    1    1    870
0    2680    7    1    2    956    870
0    2698    5    1    1    870
0    2699    7    1    2    956    870
0    2717    5    1    1    870
0    2718    7    1    2    956    870
0    2734    5    1    1    870
0    2735    7    1    2    956    870
0    2752    5    1    1    870
0    2753    7    1    2    956    870
0    2769    5    1    1    870
0    2770    7    1    2    956    870
0    2786    5    1    1    870
0    2787    7    1    2    956    870
0    2803    5    1    1    870
0    2804    7    1    2    956    870
0    359    3    1    3    917    920    923
0    1029    4    1    3    917    920    923
0    565    6    1    2    2970    2973
0    566    6    1    2    2967    2974
0    569    6    1    2    2978    2981
0    570    6    1    2    2975    2982
0    589    6    1    2    3050    3053
0    590    6    1    2    3047    3054
0    595    6    1    2    3058    3061
0    596    6    1    2    3055    3062
0    929    7    1    2    650    926
0    938    7    1    2    630    928
0    944    7    1    2    645    941
0    986    3    1    3    983    984    985
0    1014    3    1    3    1011    1012    1013
0    1616    7    1    2    442    1611
0    1625    7    1    2    456    1620
0    1634    7    1    2    463    1629
0    1643    7    1    2    479    1638
0    360    5    1    1    1029
0    567    6    1    2    565    566
0    571    6    1    2    569    570
2    579    1    576
0    591    6    1    2    589    590
0    597    6    1    2    595    596
0    614    7    1    2    576    610
0    1240    5    1    1    1075
0    1241    5    1    1    1087
0    1242    5    1    1    1099
0    1243    5    1    1    1111
0    1244    5    1    1    1123
0    1245    5    1    1    1135
0    1246    5    1    1    1147
0    1247    5    1    1    1159
0    1257    5    1    1    1075
0    1258    5    1    1    1087
0    1259    5    1    1    1099
0    1260    5    1    1    1111
0    1261    5    1    1    1123
0    1262    5    1    1    1135
0    1263    5    1    1    1147
0    1264    5    1    1    1159
0    1274    5    1    1    1075
0    1275    5    1    1    1087
0    1276    5    1    1    1099
0    1277    5    1    1    1111
0    1278    5    1    1    1123
0    1279    5    1    1    1135
0    1280    5    1    1    1147
0    1281    5    1    1    1159
0    1291    5    1    1    1075
0    1292    5    1    1    1087
0    1293    5    1    1    1099
0    1294    5    1    1    1111
0    1295    5    1    1    1123
0    1296    5    1    1    1135
0    1297    5    1    1    1147
0    1298    5    1    1    1159
0    1308    5    1    1    1075
0    1309    5    1    1    1087
0    1310    5    1    1    1099
0    1311    5    1    1    1111
0    1312    5    1    1    1123
0    1313    5    1    1    1135
0    1314    5    1    1    1147
0    1315    5    1    1    1159
0    1325    5    1    1    1075
0    1326    5    1    1    1087
0    1327    5    1    1    1099
0    1328    5    1    1    1111
0    1329    5    1    1    1123
0    1330    5    1    1    1135
0    1331    5    1    1    1147
0    1332    5    1    1    1159
0    1342    5    1    1    1075
0    1343    5    1    1    1087
0    1344    5    1    1    1099
0    1345    5    1    1    1111
0    1346    5    1    1    1123
0    1347    5    1    1    1135
0    1348    5    1    1    1147
0    1349    5    1    1    1159
0    1359    5    1    1    1075
0    1360    5    1    1    1087
0    1361    5    1    1    1099
0    1362    5    1    1    1111
0    1363    5    1    1    1123
0    1364    5    1    1    1135
0    1365    5    1    1    1147
0    1366    5    1    1    1159
0    1376    5    1    1    1168
0    1377    5    1    1    1177
0    1378    5    1    1    1186
0    1379    5    1    1    1195
0    1380    5    1    1    1204
0    1381    5    1    1    1213
0    1382    5    1    1    1222
0    1383    5    1    1    1231
0    1393    5    1    1    1168
0    1394    5    1    1    1177
0    1395    5    1    1    1186
0    1396    5    1    1    1195
0    1397    5    1    1    1204
0    1398    5    1    1    1213
0    1399    5    1    1    1222
0    1400    5    1    1    1231
0    1410    5    1    1    1168
0    1411    5    1    1    1177
0    1412    5    1    1    1186
0    1413    5    1    1    1195
0    1414    5    1    1    1204
0    1415    5    1    1    1213
0    1416    5    1    1    1222
0    1417    5    1    1    1231
0    1427    5    1    1    1168
0    1428    5    1    1    1177
0    1429    5    1    1    1186
0    1430    5    1    1    1195
0    1431    5    1    1    1204
0    1432    5    1    1    1213
0    1433    5    1    1    1222
0    1434    5    1    1    1231
0    1444    5    1    1    1168
0    1445    5    1    1    1177
0    1446    5    1    1    1186
0    1447    5    1    1    1195
0    1448    5    1    1    1204
0    1449    5    1    1    1213
0    1450    5    1    1    1222
0    1451    5    1    1    1231
0    1461    5    1    1    1168
0    1462    5    1    1    1177
0    1463    5    1    1    1186
0    1464    5    1    1    1195
0    1465    5    1    1    1204
0    1466    5    1    1    1213
0    1467    5    1    1    1222
0    1468    5    1    1    1231
0    1478    5    1    1    1168
0    1479    5    1    1    1177
0    1480    5    1    1    1186
0    1481    5    1    1    1195
0    1482    5    1    1    1204
0    1483    5    1    1    1213
0    1484    5    1    1    1222
0    1485    5    1    1    1231
0    1495    5    1    1    1168
0    1496    5    1    1    1177
0    1497    5    1    1    1186
0    1498    5    1    1    1195
0    1499    5    1    1    1204
0    1500    5    1    1    1213
0    1501    5    1    1    1222
0    1502    5    1    1    1231
2    1877    1    1874
0    1880    5    1    1    1874
0    1891    5    1    1    1866
0    1903    7    1    2    986    1901
2    1927    1    1924
0    1930    5    1    1    1924
2    1978    1    1975
0    1981    5    1    1    1975
0    1992    5    1    1    1967
2    2028    1    2025
0    2031    5    1    1    2025
0    2042    5    1    1    2017
2    2085    1    2080
0    2088    5    1    1    2080
0    2099    5    1    1    2072
0    2111    7    1    2    1014    2109
2    2137    1    2132
0    2140    5    1    1    2132
2    2190    1    2185
0    2193    5    1    1    2185
0    2204    5    1    1    2177
2    2242    1    2237
0    2245    5    1    1    2237
0    2256    5    1    1    2229
0    2320    7    1    2    2285    1862
0    2341    7    1    2    2289    1963
0    2354    7    1    2    2289    2013
0    2367    7    1    2    2289    2068
0    2383    7    1    2    2298    2173
0    2391    7    1    2    2298    2225
0    2474    5    1    1    2080
0    2475    5    1    1    2132
0    2476    5    1    1    2185
0    2477    5    1    1    2237
0    2482    7    1    5    2080    2132    2185    2237    2481
3    361    6    1    2    359    360
0    568    5    1    1    567
0    618    3    1    3    614    616    617
0    1248    7    1    2    124    1240
0    1249    7    1    2    159    1241
0    1250    7    1    2    150    1242
0    1251    7    1    2    143    1243
0    1252    7    1    2    137    1244
0    1253    7    1    2    132    1245
0    1254    7    1    2    128    1246
0    1255    7    1    2    125    1247
0    1265    7    1    2    125    1257
0    1266    7    1    2    432    1258
0    1267    7    1    2    159    1259
0    1268    7    1    2    150    1260
0    1269    7    1    2    143    1261
0    1270    7    1    2    137    1262
0    1271    7    1    2    132    1263
0    1272    7    1    2    128    1264
0    1282    7    1    2    128    1274
0    1283    7    1    2    447    1275
0    1284    7    1    2    432    1276
0    1285    7    1    2    159    1277
0    1286    7    1    2    150    1278
0    1287    7    1    2    143    1279
0    1288    7    1    2    137    1280
0    1289    7    1    2    132    1281
0    1299    7    1    2    132    1291
0    1300    7    1    2    467    1292
0    1301    7    1    2    447    1293
0    1302    7    1    2    432    1294
0    1303    7    1    2    159    1295
0    1304    7    1    2    150    1296
0    1305    7    1    2    143    1297
0    1306    7    1    2    137    1298
0    1316    7    1    2    137    1308
0    1317    7    1    2    483    1309
0    1318    7    1    2    467    1310
0    1319    7    1    2    447    1311
0    1320    7    1    2    432    1312
0    1321    7    1    2    159    1313
0    1322    7    1    2    150    1314
0    1323    7    1    2    143    1315
0    1333    7    1    2    143    1325
0    1334    7    1    2    492    1326
0    1335    7    1    2    483    1327
0    1336    7    1    2    467    1328
0    1337    7    1    2    447    1329
0    1338    7    1    2    432    1330
0    1339    7    1    2    159    1331
0    1340    7    1    2    150    1332
0    1350    7    1    2    150    1342
0    1351    7    1    2    504    1343
0    1352    7    1    2    492    1344
0    1353    7    1    2    483    1345
0    1354    7    1    2    467    1346
0    1355    7    1    2    447    1347
0    1356    7    1    2    432    1348
0    1357    7    1    2    159    1349
0    1367    7    1    2    159    1359
0    1368    7    1    2    517    1360
0    1369    7    1    2    504    1361
0    1370    7    1    2    492    1362
0    1371    7    1    2    483    1363
0    1372    7    1    2    467    1364
0    1373    7    1    2    447    1365
0    1374    7    1    2    432    1366
0    1384    7    1    2    283    1376
0    1385    7    1    2    447    1377
0    1386    7    1    2    467    1378
0    1387    7    1    2    483    1379
0    1388    7    1    2    492    1380
0    1389    7    1    2    504    1381
0    1390    7    1    2    517    1382
0    1391    7    1    2    530    1383
0    1401    7    1    2    294    1393
0    1402    7    1    2    467    1394
0    1403    7    1    2    483    1395
0    1404    7    1    2    492    1396
0    1405    7    1    2    504    1397
0    1406    7    1    2    517    1398
0    1407    7    1    2    530    1399
0    1408    7    1    2    283    1400
0    1418    7    1    2    303    1410
0    1419    7    1    2    483    1411
0    1420    7    1    2    492    1412
0    1421    7    1    2    504    1413
0    1422    7    1    2    517    1414
0    1423    7    1    2    530    1415
0    1424    7    1    2    283    1416
0    1425    7    1    2    294    1417
0    1435    7    1    2    311    1427
0    1436    7    1    2    492    1428
0    1437    7    1    2    504    1429
0    1438    7    1    2    517    1430
0    1439    7    1    2    530    1431
0    1440    7    1    2    283    1432
0    1441    7    1    2    294    1433
0    1442    7    1    2    303    1434
0    1452    7    1    2    317    1444
0    1453    7    1    2    504    1445
0    1454    7    1    2    517    1446
0    1455    7    1    2    530    1447
0    1456    7    1    2    283    1448
0    1457    7    1    2    294    1449
0    1458    7    1    2    303    1450
0    1459    7    1    2    311    1451
0    1469    7    1    2    322    1461
0    1470    7    1    2    517    1462
0    1471    7    1    2    530    1463
0    1472    7    1    2    283    1464
0    1473    7    1    2    294    1465
0    1474    7    1    2    303    1466
0    1475    7    1    2    311    1467
0    1476    7    1    2    317    1468
0    1486    7    1    2    326    1478
0    1487    7    1    2    530    1479
0    1488    7    1    2    283    1480
0    1489    7    1    2    294    1481
0    1490    7    1    2    303    1482
0    1491    7    1    2    311    1483
0    1492    7    1    2    317    1484
0    1493    7    1    2    322    1485
0    1503    7    1    2    329    1495
0    1504    7    1    2    283    1496
0    1505    7    1    2    294    1497
0    1506    7    1    2    303    1498
0    1507    7    1    2    311    1499
0    1508    7    1    2    317    1500
0    1509    7    1    2    322    1501
0    1510    7    1    2    326    1502
0    2483    7    1    5    2474    2475    2476    2477    2478
2    600    1    597
0    661    7    1    2    568    660
0    669    7    1    2    597    665
0    679    7    1    2    591    678
0    1256    4    1    8    1248    1249    1250    1251    1252    1253    1254    1255
0    1273    4    1    8    1265    1266    1267    1268    1269    1270    1271    1272
0    1290    4    1    8    1282    1283    1284    1285    1286    1287    1288    1289
0    1307    4    1    8    1299    1300    1301    1302    1303    1304    1305    1306
0    1324    4    1    8    1316    1317    1318    1319    1320    1321    1322    1323
0    1341    4    1    8    1333    1334    1335    1336    1337    1338    1339    1340
0    1358    4    1    8    1350    1351    1352    1353    1354    1355    1356    1357
0    1375    4    1    8    1367    1368    1369    1370    1371    1372    1373    1374
0    1392    4    1    8    1384    1385    1386    1387    1388    1389    1390    1391
0    1409    4    1    8    1401    1402    1403    1404    1405    1406    1407    1408
0    1426    4    1    8    1418    1419    1420    1421    1422    1423    1424    1425
0    1443    4    1    8    1435    1436    1437    1438    1439    1440    1441    1442
0    1460    4    1    8    1452    1453    1454    1455    1456    1457    1458    1459
0    1477    4    1    8    1469    1470    1471    1472    1473    1474    1475    1476
0    1494    4    1    8    1486    1487    1488    1489    1490    1491    1492    1493
0    1511    4    1    8    1503    1504    1505    1506    1507    1508    1509    1510
0    1652    7    1    2    618    1647
0    1883    7    1    3    169    1862    1877
0    1886    7    1    3    179    1862    1880
0    1889    7    1    3    190    1866    1880
0    1890    7    1    3    200    1866    1877
0    1912    3    1    3    1903    1906    1909
0    1916    4    1    3    1903    1906    1909
0    1984    7    1    3    169    1963    1978
0    1987    7    1    3    179    1963    1981
0    1990    7    1    3    190    1967    1981
0    1991    7    1    3    200    1967    1978
0    2034    7    1    3    169    2013    2028
0    2037    7    1    3    179    2013    2031
0    2040    7    1    3    190    2017    2031
0    2041    7    1    3    200    2017    2028
0    2091    7    1    3    169    2068    2085
0    2094    7    1    3    179    2068    2088
0    2097    7    1    3    190    2072    2088
0    2098    7    1    3    200    2072    2085
0    2120    3    1    3    2111    2114    2117
0    2124    4    1    3    2111    2114    2117
0    2196    7    1    3    169    2173    2190
0    2199    7    1    3    179    2173    2193
0    2202    7    1    3    190    2177    2193
0    2203    7    1    3    200    2177    2190
0    2248    7    1    3    169    2225    2242
0    2251    7    1    3    179    2225    2245
0    2254    7    1    3    190    2229    2245
0    2255    7    1    3    200    2229    2242
0    2484    3    1    2    2482    2483
2    2991    1    571
2    2994    1    579
2    2999    1    571
2    3002    1    579
2    3063    1    591
2    3071    1    591
2    3124    1    2320
2    3134    1    2320
2    3158    1    2341
2    3166    1    2341
2    3174    1    2354
2    3182    1    2354
2    3190    1    2367
2    3200    1    2367
2    3224    1    2383
2    3232    1    2383
2    3240    1    2391
2    3248    1    2391
0    663    4    1    2    661    662
0    673    3    1    3    669    671    672
0    681    4    1    2    679    680
0    1536    7    1    2    1256    1533
0    1537    7    1    2    1392    1534
0    1582    7    1    2    1273    1581
0    1583    7    1    2    1409    1512
0    1586    7    1    2    1290    1585
0    1587    7    1    2    1426    1512
0    1590    7    1    2    1307    1589
0    1591    7    1    2    1443    1512
0    1594    7    1    2    1324    1593
0    1595    7    1    2    1460    1512
0    1598    7    1    2    1341    1597
0    1599    7    1    2    1477    1512
0    1602    7    1    2    1358    1601
0    1603    7    1    2    1494    1512
0    1606    7    1    2    1375    1605
0    1607    7    1    2    1511    1512
0    1894    3    1    3    1889    1890    1891
0    1997    3    1    3    1990    1991    1992
0    2047    3    1    3    2040    2041    2042
0    2102    3    1    3    2097    2098    2099
0    2209    3    1    3    2202    2203    2204
0    2261    3    1    3    2254    2255    2256
0    2489    7    1    2    2484    2488
0    3005    5    1    1    2999
0    3006    5    1    1    3002
0    3077    5    1    1    3071
0    3069    5    1    1    3063
0    2997    5    1    1    2991
0    2998    5    1    1    2994
0    689    7    1    2    681    683
0    700    7    1    2    663    694
0    1539    3    1    3    1536    1537    1538
0    1584    3    1    2    1582    1583
0    1588    3    1    2    1586    1587
0    1592    3    1    2    1590    1591
0    1596    3    1    2    1594    1595
0    1600    3    1    2    1598    1599
0    1604    3    1    2    1602    1603
0    1608    3    1    2    1606    1607
0    1661    7    1    2    673    1656
0    1892    3    1    2    1883    1886
0    1893    4    1    2    1883    1886
0    1933    7    1    3    169    1912    1927
0    1936    7    1    3    179    1912    1930
0    1939    7    1    3    190    1916    1930
0    1940    7    1    3    200    1916    1927
0    1941    5    1    1    1916
0    1993    3    1    2    1984    1987
0    1996    4    1    2    1984    1987
0    2043    3    1    2    2034    2037
0    2046    4    1    2    2034    2037
0    2100    3    1    2    2091    2094
0    2101    4    1    2    2091    2094
0    2143    7    1    3    169    2120    2137
0    2146    7    1    3    179    2120    2140
0    2149    7    1    3    190    2124    2140
0    2150    7    1    3    200    2124    2137
0    2151    5    1    1    2124
0    2205    3    1    2    2196    2199
0    2208    4    1    2    2196    2199
0    2257    3    1    2    2248    2251
0    2260    4    1    2    2248    2251
0    3138    5    1    1    3134
0    2328    7    1    2    2285    1912
0    3162    5    1    1    3158
0    3170    5    1    1    3166
0    3178    5    1    1    3174
0    3186    5    1    1    3182
0    3204    5    1    1    3200
0    2375    7    1    2    2298    2120
0    3236    5    1    1    3232
0    3244    5    1    1    3240
0    3252    5    1    1    3248
0    3228    5    1    1    3224
2    3066    1    600
2    3074    1    600
0    3128    5    1    1    3124
0    3194    5    1    1    3190
0    619    6    1    2    2994    2997
0    620    6    1    2    2991    2998
0    582    6    1    2    3002    3005
0    583    6    1    2    2999    3006
0    692    3    1    3    689    690    691
0    703    3    1    3    700    701    702
0    1612    7    1    2    1539    1609
0    1621    7    1    2    1584    1618
0    1630    7    1    2    1588    1627
0    1639    7    1    2    1592    1636
0    1648    7    1    2    1596    1645
0    1657    7    1    2    1600    1654
0    1666    7    1    2    1604    1663
0    1675    7    1    2    1608    1672
0    1895    7    1    2    1893    1894
0    1946    3    1    3    1939    1940    1941
0    1998    7    1    2    1996    1997
0    2048    7    1    2    2046    2047
0    2103    7    1    2    2101    2102
0    2156    3    1    3    2149    2150    2151
0    2210    7    1    2    2208    2209
0    2262    7    1    2    2260    2261
0    2271    5    1    1    1892
0    2311    5    1    1    2100
0    356    6    1    2    619    620
0    357    6    1    2    582    583
0    603    6    1    2    3074    3077
0    3078    5    1    1    3074
0    606    6    1    2    3066    3069
0    3070    5    1    1    3066
0    1670    7    1    2    703    1665
0    1679    7    1    2    692    1674
0    1942    3    1    2    1933    1936
0    1945    4    1    2    1933    1936
0    2152    3    1    2    2143    2146
0    2155    4    1    2    2143    2146
0    2445    7    1    2    1993    2293
0    2448    7    1    2    2043    2293
0    2455    7    1    2    2205    2302
0    2458    7    1    2    2257    2302
2    3142    1    2328
2    3150    1    2328
2    3208    1    2375
2    3216    1    2375
3    358    6    1    2    356    357
0    604    6    1    2    3071    3078
0    607    6    1    2    3063    3070
0    1947    7    1    2    1945    1946
0    2157    7    1    2    2155    2156
2    2317    1    1895
2    2338    1    1998
2    2351    1    2048
2    2364    1    2103
2    2380    1    2210
2    2388    1    2262
0    605    6    1    2    603    604
0    608    6    1    2    606    607
0    2272    6    1    2    1895    1942
0    2312    6    1    2    2103    2152
0    3146    5    1    1    3142
0    3154    5    1    1    3150
0    3220    5    1    1    3216
0    3212    5    1    1    3208
0    2444    7    1    2    1942    2288
2    2451    1    2448
0    2454    7    1    2    2152    2293
2    2461    1    2458
0    2530    5    1    1    2445
2    3323    1    2458
0    349    5    1    1    605
0    350    5    1    1    608
0    2265    7    1    4    1895    1947    1998    2048
0    2273    6    1    3    1895    1947    1993
0    2274    6    1    4    2043    1947    1998    1895
0    2309    7    1    4    2103    2157    2210    2262
0    2313    6    1    3    2103    2157    2205
0    2314    6    1    4    2257    2157    2210    2103
2    2325    1    1947
2    2372    1    2157
0    2523    5    1    1    2444
0    2533    5    1    1    2454
2    3121    1    2317
2    3131    1    2317
2    3155    1    2338
2    3163    1    2338
2    3171    1    2351
2    3179    1    2351
2    3187    1    2364
2    3197    1    2364
2    3221    1    2380
2    3229    1    2380
2    3237    1    2388
2    3245    1    2388
3    351    6    1    2    349    350
0    2275    6    1    4    2271    2272    2273    2274
0    2315    6    1    4    2311    2312    2313    2314
0    3329    5    1    1    3323
3    372    7    1    2    2309    2265
0    2324    6    1    2    3131    3138
0    2350    6    1    2    3163    3170
0    2363    6    1    2    3179    3186
0    2371    6    1    2    3197    3204
0    2387    6    1    2    3229    3236
0    2400    6    1    2    3245    3252
2    2268    1    2265
0    3137    5    1    1    3131
0    3161    5    1    1    3155
0    2345    6    1    2    3155    3162
0    3169    5    1    1    3163
0    3177    5    1    1    3171
0    2358    6    1    2    3171    3178
0    3185    5    1    1    3179
0    3203    5    1    1    3197
0    3235    5    1    1    3229
0    3243    5    1    1    3237
0    2395    6    1    2    3237    3244
0    3251    5    1    1    3245
0    3227    5    1    1    3221
0    2432    6    1    2    3221    3228
0    2490    7    1    2    2309    2485
0    3127    5    1    1    3121
0    3130    6    1    2    3121    3128
2    3139    1    2325
2    3147    1    2325
0    3193    5    1    1    3187
0    3196    6    1    2    3187    3194
2    3205    1    2372
2    3213    1    2372
0    2307    6    1    2    2265    2315
0    2308    5    1    1    2275
0    2323    6    1    2    3134    3137
0    2349    6    1    2    3166    3169
0    2362    6    1    2    3182    3185
0    2370    6    1    2    3200    3203
0    2386    6    1    2    3232    3235
0    2399    6    1    2    3248    3251
0    2344    6    1    2    3158    3161
0    2357    6    1    2    3174    3177
0    2394    6    1    2    3240    3243
0    2431    6    1    2    3224    3227
0    2464    7    1    2    2315    2302
0    2491    3    1    2    2489    2490
0    3129    6    1    2    3124    3127
0    3195    6    1    2    3190    3193
0    368    7    1    2    2307    2308
0    1615    6    1    2    2323    2324
0    2337    6    1    2    3147    3154
0    1633    6    1    2    2349    2350
0    1642    6    1    2    2362    2363
0    1651    6    1    2    2370    2371
0    2379    6    1    2    3213    3220
0    1669    6    1    2    2386    2387
0    1678    6    1    2    2399    2400
0    3145    5    1    1    3139
0    2332    6    1    2    3139    3146
0    3153    5    1    1    3147
0    2346    6    1    2    2344    2345
0    2359    6    1    2    2357    2358
0    3219    5    1    1    3213
0    2396    6    1    2    2394    2395
0    3211    5    1    1    3205
0    2425    6    1    2    3205    3212
0    2433    6    1    2    2431    2432
0    3272    6    1    2    3129    3130
0    3308    6    1    2    3195    3196
3    369    5    1    1    368
0    1613    5    1    1    1615
0    2336    6    1    2    3150    3153
0    1631    5    1    1    1633
0    1640    5    1    1    1642
0    1649    5    1    1    1651
0    2378    6    1    2    3216    3219
0    1667    5    1    1    1669
0    1676    5    1    1    1678
0    2331    6    1    2    3142    3145
0    2424    6    1    2    3208    3211
2    2467    1    2464
2    2495    1    2491
2    3295    1    2464
0    3374    7    1    2    330    2491
0    1614    7    1    2    1613    1610
0    1624    6    1    2    2336    2337
0    1632    7    1    2    1631    1628
0    1641    7    1    2    1640    1637
0    1650    7    1    2    1649    1646
0    1660    6    1    2    2378    2379
0    1668    7    1    2    1667    1664
0    1677    7    1    2    1676    1673
0    2333    6    1    2    2331    2332
2    2406    1    2346
2    2409    1    2346
2    2415    1    2359
2    2419    1    2359
0    2426    6    1    2    2424    2425
2    2439    1    2396
0    2518    7    1    2    2433    2461
0    3276    5    1    1    3272
0    3312    5    1    1    3308
0    2612    7    1    2    330    2396
2    3326    1    2433
0    1617    4    1    3    1612    1614    1616
0    1622    5    1    1    1624
0    1635    4    1    3    1630    1632    1634
0    1644    4    1    3    1639    1641    1643
0    1653    4    1    3    1648    1650    1652
0    1658    5    1    1    1660
0    1671    4    1    3    1666    1668    1670
0    1680    4    1    3    1675    1677    1679
0    2500    7    1    2    2467    2268
0    2505    7    1    2    2495    2268
0    2519    3    1    2    2455    2518
0    3378    5    1    1    3374
0    2642    5    1    1    2467
2    2645    1    2467
0    3301    5    1    1    3295
0    1623    7    1    2    1622    1619
0    1659    7    1    2    1658    1655
2    2401    1    2333
0    2501    3    1    2    2275    2500
0    2511    7    1    3    2495    2419    2409
0    2512    7    1    2    2495    2415
0    2513    7    1    3    2439    2433    2426
0    2514    7    1    2    2439    2433
0    2517    7    1    2    2467    2415
0    2531    6    1    2    2409    2451
0    2532    6    1    3    2409    2419    2467
0    2534    6    1    2    2426    2455
0    2535    6    1    3    2426    2433    2461
0    2607    6    1    2    3326    3329
0    3330    5    1    1    3326
0    2643    7    1    3    330    2491    2642
0    2687    7    1    2    1617    2680
0    2725    7    1    2    1635    2718
0    2742    7    1    2    1644    2735
0    2760    7    1    2    1653    2753
0    2794    7    1    2    1671    2787
0    2811    7    1    2    1680    2804
2    3280    1    2333
2    3290    1    2409
2    3298    1    2415
2    3316    1    2426
2    3406    1    2612
2    3414    1    2612
0    3422    7    1    2    2439    2439
0    1626    4    1    3    1621    1623    1625
0    1662    4    1    3    1657    1659    1661
0    2567    7    1    2    330    2512
0    2589    7    1    2    330    2513
0    2608    6    1    2    3323    3330
2    2654    1    2519
2    3253    1    2505
0    3277    6    1    3    2530    2531    2532
0    3287    3    1    2    2448    2517
0    3305    6    1    3    2533    2534    2535
2    3313    1    2519
0    3350    7    1    2    330    2511
0    932    3    1    2    2643    2645
0    2508    7    1    4    2495    2401    2409    2419
0    2524    6    1    2    2401    2445
0    2525    6    1    3    2401    2406    2451
0    2526    6    1    4    2401    2406    2419    2467
0    3294    5    1    1    3290
0    2609    6    1    2    2607    2608
0    3410    5    1    1    3406
0    3418    5    1    1    3414
0    2624    6    1    2    3422    3425
0    3426    5    1    1    3422
2    2629    1    2501
0    2647    4    1    2    2643    2645
0    2706    7    1    2    1626    2699
0    2777    7    1    2    1662    2770
2    3264    1    2501
0    3284    5    1    1    3280
0    3302    5    1    1    3298
0    3303    6    1    2    3298    3301
0    3320    5    1    1    3316
0    3398    7    1    2    330    2514
0    2657    5    1    1    2654
0    398    7    1    2    2519    2654
0    933    7    1    2    932    927
0    2527    6    1    4    2523    2524    2525    2526
0    3259    5    1    1    3253
0    3354    5    1    1    3350
0    3293    5    1    1    3287
0    2563    6    1    2    3287    3294
0    3311    5    1    1    3305
0    2585    6    1    2    3305    3312
0    2625    6    1    2    3419    3426
0    3283    5    1    1    3277
0    3286    6    1    2    3277    3284
0    3304    6    1    2    3295    3302
0    3319    5    1    1    3313
0    3322    6    1    2    3313    3320
2    3358    1    2567
2    3366    1    2567
2    3382    1    2589
2    3390    1    2589
0    397    7    1    3    330    2514    2657
0    2544    7    1    2    330    2508
0    2562    6    1    2    3290    3293
0    2584    6    1    2    3308    3311
0    3402    5    1    1    3398
0    2626    6    1    2    2624    2625
0    2632    5    1    1    2629
0    2634    7    1    2    2501    2629
2    2650    1    2647
0    3268    5    1    1    3264
2    3256    1    2508
0    3285    6    1    2    3280    3283
0    3321    6    1    2    3316    3319
0    3371    6    1    2    3303    3304
2    3403    1    2609
2    3411    1    2609
0    362    3    1    3    929    933    938
0    1030    4    1    3    929    933    938
3    399    3    1    2    397    398
0    2564    6    1    2    2562    2563
0    3362    5    1    1    3358
0    3370    5    1    1    3366
0    2586    6    1    2    2584    2585
0    3386    5    1    1    3382
0    3394    5    1    1    3390
0    2633    7    1    3    330    2505    2632
2    3261    1    2527
2    3269    1    2527
0    3347    6    1    2    3285    3286
0    3395    6    1    2    3321    3322
0    363    5    1    1    1030
0    2536    6    1    2    3256    3259
0    3260    5    1    1    3256
0    3377    5    1    1    3371
0    2580    6    1    2    3371    3378
0    3409    5    1    1    3403
0    2616    6    1    2    3403    3410
0    3417    5    1    1    3411
0    2622    6    1    2    3411    3418
0    2635    4    1    2    2633    2634
0    2805    7    1    2    2626    2802
0    2808    7    1    2    2626    2803
2    3334    1    2544
2    3342    1    2544
2    3454    1    2650
3    364    7    1    2    362    363
0    2537    6    1    2    3253    3260
0    3275    5    1    1    3269
0    2540    6    1    2    3269    3276
0    3353    5    1    1    3347
0    2557    6    1    2    3347    3354
0    2579    6    1    2    3374    3377
0    3401    5    1    1    3395
0    2602    6    1    2    3395    3402
0    2615    6    1    2    3406    3409
0    2621    6    1    2    3414    3417
0    3267    5    1    1    3261
0    3112    6    1    2    3261    3268
2    3355    1    2564
2    3363    1    2564
2    3379    1    2586
2    3387    1    2586
0    2538    6    1    2    2536    2537
0    2539    6    1    2    3272    3275
0    3338    5    1    1    3334
0    3346    5    1    1    3342
0    2556    6    1    2    3350    3353
0    2581    6    1    2    2579    2580
0    2601    6    1    2    3398    3401
0    2617    6    1    2    2615    2616
0    2623    6    1    2    2621    2622
2    2638    1    2635
0    3458    5    1    1    3454
0    2814    3    1    3    2805    2808    2811
0    2816    4    1    3    2805    2808    2811
0    3111    6    1    2    3264    3267
0    2541    6    1    2    2539    2540
0    2558    6    1    2    2556    2557
0    3361    5    1    1    3355
0    2571    6    1    2    3355    3362
0    3369    5    1    1    3363
0    2577    6    1    2    3363    3370
0    3385    5    1    1    3379
0    2593    6    1    2    3379    3386
0    3393    5    1    1    3387
0    2598    6    1    2    3387    3394
0    2603    6    1    2    2601    2602
0    3113    6    1    2    3111    3112
0    3116    7    1    2    330    2538
0    3451    5    1    1    2623
0    395    5    1    1    2816
0    2570    6    1    2    3358    3361
0    2576    6    1    2    3366    3369
0    2592    6    1    2    3382    3385
0    2597    6    1    2    3390    3393
0    2736    7    1    2    2581    2733
0    2739    7    1    2    2581    2734
0    2788    7    1    2    2617    2785
2    3438    1    2638
0    3446    7    1    2    2617    2647
2    3459    1    2814
3    396    7    1    2    2814    395
0    3119    5    1    1    3113
0    3120    5    1    1    3116
0    2572    6    1    2    2570    2571
0    2578    6    1    2    2576    2577
0    2594    6    1    2    2592    2593
0    2599    6    1    2    2597    2598
0    2677    6    1    2    3451    3458
0    3457    5    1    1    3451
0    2700    7    1    2    2558    2697
0    2771    7    1    2    2603    2768
2    3331    1    2541
2    3339    1    2541
2    3427    1    2558
2    3443    1    2603
0    954    6    1    2    3116    3119
0    955    6    1    2    3113    3120
0    2600    5    1    1    2599
0    3442    5    1    1    3438
0    3450    5    1    1    3446
0    2676    6    1    2    3454    3457
0    2745    3    1    3    2736    2739    2742
0    2748    4    1    3    2736    2739    2742
0    3465    5    1    1    3459
0    3435    5    1    1    2578
0    950    6    1    2    954    955
0    3337    5    1    1    3331
0    2548    6    1    2    3331    3338
0    3345    5    1    1    3339
0    2553    6    1    2    3339    3346
0    2661    4    1    2    2600    2650
0    2662    7    1    4    2617    2603    2594    2650
0    3433    5    1    1    3427
0    3449    5    1    1    3443
0    2672    6    1    2    3443    3450
0    2674    6    1    2    2676    2677
0    2719    7    1    2    2572    2716
0    2754    7    1    2    2594    2751
0    3430    7    1    2    2572    2635
0    383    5    1    1    2748
0    951    7    1    2    950    943
0    2547    6    1    2    3334    3337
0    2552    6    1    2    3342    3345
0    2663    3    1    2    2661    2662
0    2670    6    1    2    3435    3442
0    3441    5    1    1    3435
0    2671    6    1    2    3446    3449
0    2675    5    1    1    2674
2    3491    1    2745
2    3499    1    2745
3    384    7    1    2    2745    383
0    2549    6    1    2    2547    2548
0    2554    6    1    2    2552    2553
0    2664    6    1    2    3430    3433
0    3434    5    1    1    3430
0    2669    6    1    2    3438    3441
0    2673    6    1    2    2671    2672
0    2757    7    1    2    2663    2752
0    2791    7    1    2    2675    2786
0    365    3    1    3    944    947    951
0    1031    4    1    3    944    947    951
0    2555    5    1    1    2554
0    2665    6    1    2    3427    3434
0    2667    6    1    2    2669    2670
0    2774    7    1    2    2673    2769
0    3497    5    1    1    3491
0    3505    5    1    1    3499
0    366    5    1    1    1031
0    2658    4    1    2    2555    2638
0    2659    7    1    4    2572    2558    2549    2638
0    2666    6    1    2    2664    2665
0    2668    5    1    1    2667
0    2681    7    1    2    2549    2678
0    2763    3    1    3    2754    2757    2760
0    2765    4    1    3    2754    2757    2760
0    2797    3    1    3    2788    2791    2794
0    2799    4    1    3    2788    2791    2794
3    367    7    1    2    365    366
0    2660    3    1    2    2658    2659
0    2703    7    1    2    2666    2698
0    2722    7    1    2    2668    2717
0    2780    3    1    3    2771    2774    2777
0    2782    4    1    3    2771    2774    2777
0    386    5    1    1    2765
0    392    5    1    1    2799
0    2684    7    1    2    2660    2679
2    3462    1    2797
2    3470    1    2763
3    387    7    1    2    2763    386
0    389    5    1    1    2782
3    393    7    1    2    2797    392
0    2709    3    1    3    2700    2703    2706
0    2713    4    1    3    2700    2703    2706
0    2728    3    1    3    2719    2722    2725
0    2730    4    1    3    2719    2722    2725
0    2922    7    1    4    2816    2799    2782    2765
2    3467    1    2780
3    390    7    1    2    2780    389
0    2690    3    1    3    2681    2684    2687
0    2694    4    1    3    2681    2684    2687
0    2821    6    1    2    3462    3465
0    3466    5    1    1    3462
0    3474    5    1    1    3470
3    378    7    1    2    2709    2709
0    380    5    1    1    2730
0    2822    6    1    2    3459    3466
0    3473    5    1    1    3467
0    2827    6    1    2    3467    3474
2    2839    1    2728
0    2883    7    1    2    2709    2871
2    3507    1    2709
3    375    7    1    2    2690    2690
3    381    7    1    2    2728    380
0    2823    6    1    2    2821    2822
0    2826    6    1    2    3470    3473
0    2880    7    1    2    2871    2690
0    2925    7    1    4    2748    2730    2713    2694
0    2928    7    1    3    2713    2694    2874
2    3510    1    2690
0    2828    6    1    2    2826    2827
2    3494    1    2839
2    3502    1    2839
0    3513    5    1    1    3507
2    3544    1    2883
2    3552    1    2883
0    406    7    1    2    2922    2925
0    2929    7    1    2    2922    2925
2    3475    1    2823
2    3483    1    2823
0    3514    5    1    1    3510
0    3515    6    1    2    3510    3513
2    3541    1    2880
2    3549    1    2880
3    407    5    1    1    406
0    2930    4    1    2    2928    2929
0    2842    6    1    2    3494    3497
0    3498    5    1    1    3494
0    2852    6    1    2    3502    3505
0    3506    5    1    1    3502
0    3548    5    1    1    3544
0    3556    5    1    1    3552
2    3478    1    2828
2    3486    1    2828
0    3516    6    1    2    3507    3514
0    408    7    1    2    213    2930
0    3481    5    1    1    3475
0    3489    5    1    1    3483
0    2843    6    1    2    3491    3498
0    2853    6    1    2    3499    3506
0    3547    5    1    1    3541
0    2887    6    1    2    3541    3548
0    2896    6    1    2    3549    3556
0    3555    5    1    1    3549
0    3520    6    1    2    3515    3516
3    409    5    1    1    408
0    2831    6    1    2    3478    3481
0    3482    5    1    1    3478
0    2836    6    1    2    3486    3489
0    3490    5    1    1    3486
0    2844    6    1    2    2842    2843
0    2848    6    1    2    2852    2853
0    2886    6    1    2    3544    3547
0    2895    6    1    2    3552    3555
0    2832    6    1    2    3475    3482
0    2837    6    1    2    3483    3490
0    2849    5    1    1    2848
0    3524    5    1    1    3520
0    2888    6    1    2    2886    2887
0    2891    6    1    2    2895    2896
0    2833    6    1    2    2831    2832
0    2838    6    1    2    2836    2837
0    2892    5    1    1    2891
2    3517    1    2844
0    2906    7    1    3    2844    2888    2900
0    2908    7    1    3    2849    2888    2903
0    2913    5    1    1    2838
0    3523    5    1    1    3517
0    2855    6    1    2    3517    3524
0    2907    7    1    3    2844    2892    2903
0    2909    7    1    3    2849    2892    2900
2    3525    1    2833
2    3533    1    2833
0    2854    6    1    2    3520    3523
0    2910    3    1    4    2906    2907    2908    2909
2    3560    1    2913
2    3568    1    2913
0    2856    6    1    2    2854    2855
0    3539    5    1    1    3533
0    3531    5    1    1    3525
0    3572    5    1    1    3568
0    3564    5    1    1    3560
2    3557    1    2910
2    3565    1    2910
2    3528    1    2856
2    3536    1    2856
0    2921    6    1    2    3557    3564
0    2917    6    1    2    3565    3572
0    3571    5    1    1    3565
0    3563    5    1    1    3557
0    2863    6    1    2    3528    3531
0    2859    6    1    2    3536    3539
0    2920    6    1    2    3560    3563
0    2916    6    1    2    3568    3571
0    3540    5    1    1    3536
0    3532    5    1    1    3528
0    2864    6    1    2    3525    3532
0    2860    6    1    2    3533    3540
0    403    6    1    2    2920    2921
0    404    6    1    2    2916    2917
0    400    6    1    2    2863    2864
0    401    6    1    2    2859    2860
3    405    7    1    2    403    404
3    402    6    1    2    400    401
