1    76    0    1    0
1    40    0    1    0
1    56    0    1    0
1    11    0    1    0
1    34    0    1    0
1    30    0    1    0
1    69    0    1    0
1    73    0    1    0
1    108    0    1    0
1    24    0    1    0
1    92    0    1    0
1    8    0    1    0
1    17    0    1    0
1    21    0    1    0
1    82    0    1    0
1    95    0    1    0
1    4    0    1    0
1    27    0    1    0
1    14    0    1    0
1    66    0    1    0
1    89    0    1    0
1    86    0    1    0
1    79    0    1    0
1    105    0    1    0
1    53    0    1    0
1    60    0    1    0
1    37    0    1    0
1    47    0    1    0
1    102    0    1    0
1    112    0    1    0
1    50    0    1    0
1    63    0    1    0
1    99    0    1    0
1    1    0    1    0
1    43    0    1    0
1    115    0    1    0
0    118    5    1    1    1
0    119    5    2    1    4
0    122    5    1    1    11
0    123    5    2    1    17
0    126    5    1    1    24
0    127    5    2    1    30
0    130    5    1    1    37
0    131    5    2    1    43
0    134    5    1    1    50
0    135    5    2    1    56
0    138    5    1    1    63
0    139    5    2    1    69
0    142    5    1    1    76
0    143    5    2    1    82
0    146    5    1    1    89
0    147    5    2    1    95
0    150    5    1    1    102
0    151    5    2    1    108
0    154    6    2    2    118    4
0    157    4    1    2    8    119
0    158    4    1    2    14    119
0    159    6    2    2    122    17
0    162    6    2    2    126    30
0    165    6    2    2    130    43
0    168    6    2    2    134    56
0    171    6    2    2    138    69
0    174    6    2    2    142    82
0    177    6    2    2    146    95
0    180    6    2    2    150    108
0    183    4    1    2    21    123
0    184    4    1    2    27    123
0    185    4    1    2    34    127
0    186    4    1    2    40    127
0    187    4    1    2    47    131
0    188    4    1    2    53    131
0    189    4    1    2    60    135
0    190    4    1    2    66    135
0    191    4    1    2    73    139
0    192    4    1    2    79    139
0    193    4    1    2    86    143
0    194    4    1    2    92    143
0    195    4    1    2    99    147
0    196    4    1    2    105    147
0    197    4    1    2    112    151
0    198    4    1    2    115    151
0    199    7    3    9    154    159    162    165    168    171    174    177    180
0    203    5    9    1    199
0    213    5    9    1    199
3    223    5    0    1    199
0    224    2    2    2    203    154
0    227    2    2    2    203    159
0    230    2    2    2    203    162
0    233    2    2    2    203    165
0    236    2    2    2    203    168
0    239    2    2    2    203    171
0    242    6    1    2    1    213
0    243    2    2    2    203    174
0    246    6    1    2    213    11
0    247    2    2    2    203    177
0    250    6    1    2    213    24
0    251    2    2    2    203    180
0    254    6    1    2    213    37
0    255    6    1    2    213    50
0    256    6    1    2    213    63
0    257    6    1    2    213    76
0    258    6    1    2    213    89
0    259    6    1    2    213    102
0    260    6    2    2    224    157
0    263    6    1    2    224    158
0    264    6    2    2    227    183
0    267    6    2    2    230    185
0    270    6    2    2    233    187
0    273    6    2    2    236    189
0    276    6    2    2    239    191
0    279    6    2    2    243    193
0    282    6    2    2    247    195
0    285    6    2    2    251    197
0    288    6    1    2    227    184
0    289    6    1    2    230    186
0    290    6    1    2    233    188
0    291    6    1    2    236    190
0    292    6    1    2    239    192
0    293    6    1    2    243    194
0    294    6    1    2    247    196
0    295    6    1    2    251    198
0    296    7    3    9    260    264    267    270    273    276    279    282    285
0    300    5    1    1    263
0    301    5    1    1    288
0    302    5    1    1    289
0    303    5    1    1    290
0    304    5    1    1    291
0    305    5    1    1    292
0    306    5    1    1    293
0    307    5    1    1    294
0    308    5    1    1    295
0    309    5    9    1    296
0    319    5    9    1    296
3    329    5    0    1    296
0    330    2    1    2    309    260
0    331    2    1    2    309    264
0    332    2    1    2    309    267
0    333    2    1    2    309    270
0    334    6    1    2    8    319
0    335    2    1    2    309    273
0    336    6    1    2    319    21
0    337    2    1    2    309    276
0    338    6    1    2    319    34
0    339    2    1    2    309    279
0    340    6    1    2    319    47
0    341    2    1    2    309    282
0    342    6    1    2    319    60
0    343    2    1    2    309    285
0    344    6    1    2    319    73
0    345    6    1    2    319    86
0    346    6    1    2    319    99
0    347    6    1    2    319    112
0    348    6    1    2    330    300
0    349    6    1    2    331    301
0    350    6    1    2    332    302
0    351    6    1    2    333    303
0    352    6    1    2    335    304
0    353    6    1    2    337    305
0    354    6    1    2    339    306
0    355    6    1    2    341    307
0    356    6    1    2    343    308
0    357    7    2    9    348    349    350    351    352    353    354    355    356
0    360    5    9    1    357
3    370    5    0    1    357
0    371    6    1    2    14    360
0    372    6    1    2    360    27
0    373    6    1    2    360    40
0    374    6    1    2    360    53
0    375    6    1    2    360    66
0    376    6    1    2    360    79
0    377    6    1    2    360    92
0    378    6    1    2    360    105
0    379    6    1    2    360    115
0    380    6    1    4    4    242    334    371
0    381    6    4    4    246    336    372    17
0    386    6    6    4    250    338    373    30
0    393    6    5    4    254    340    374    43
0    399    6    4    4    255    342    375    56
0    404    6    2    4    256    344    376    69
0    407    6    3    4    257    345    377    82
0    411    6    2    4    258    346    378    95
0    414    6    1    4    259    347    379    108
0    415    5    1    1    380
0    416    7    1    8    381    386    393    399    404    407    411    414
0    417    5    1    1    393
0    418    5    1    1    404
0    419    5    1    1    407
0    420    5    1    1    411
3    421    4    0    2    415    416
0    422    6    2    2    386    417
0    425    6    2    4    386    393    418    399
0    428    6    1    3    399    393    419
0    429    6    1    4    386    393    407    420
3    430    6    0    4    381    386    422    399
3    431    6    0    4    381    386    425    428
3    432    6    0    4    381    422    425    429
