1    274    0    1    0
1    266    0    1    0
1    2446    0    2    0
1    191    0    1    0
1    44    0    2    0
1    265    0    1    0
1    74    0    2    0
1    268    0    1    0
1    34    0    2    0
1    567    0    2    0
1    24    0    2    0
1    85    0    2    0
1    126    0    2    0
1    88    0    2    0
1    8    0    2    0
1    1981    0    2    0
1    264    0    1    0
1    118    0    2    0
1    1956    0    2    0
1    64    0    2    0
1    20    0    2    0
1    271    0    1    0
1    184    0    1    0
1    95    0    2    0
1    213    0    1    0
1    27    0    2    0
1    68    0    2    0
1    51    0    2    0
1    75    0    2    0
1    131    0    2    0
1    273    0    1    0
1    214    0    1    0
1    1991    0    2    0
1    203    0    1    0
1    2451    0    2    0
1    181    0    1    0
1    483    0    2    0
1    16    0    2    0
1    240    0    1    0
1    81    0    2    0
1    2100    0    2    0
1    207    0    1    0
1    205    0    1    0
1    2090    0    2    0
1    91    0    2    0
1    267    0    1    0
1    52    0    2    0
1    26    0    2    0
1    102    0    2    0
1    112    0    2    0
1    1348    0    2    0
1    50    0    2    0
1    1    0    2    0
1    136    0    2    0
1    23    0    2    0
1    278    0    1    0
1    256    0    1    0
1    860    0    2    0
1    101    0    2    0
1    2427    0    2    0
1    56    0    2    0
1    62    0    2    0
1    1384    0    2    0
1    868    0    2    0
1    117    0    2    0
1    108    0    2    0
1    140    0    2    0
1    3    0    2    0
1    22    0    2    0
1    48    0    2    0
1    104    0    2    0
1    246    0    1    0
1    138    0    2    0
1    125    0    2    0
1    257    0    1    0
1    183    0    1    0
1    21    0    2    0
1    137    0    2    0
1    96    0    2    0
1    279    0    1    0
1    35    0    2    0
1    77    0    2    0
1    87    0    2    0
1    113    0    2    0
1    2443    0    2    0
1    180    0    1    0
1    263    0    1    0
1    57    0    2    0
1    103    0    2    0
1    86    0    2    0
1    195    0    1    0
1    245    0    1    0
1    243    0    1    0
1    141    0    2    0
1    80    0    2    0
1    94    0    2    0
1    1083    0    2    0
1    105    0    2    0
1    248    0    1    0
1    1966    0    2    0
1    142    0    2    0
1    33    0    2    0
1    2438    0    2    0
1    67    0    2    0
1    128    0    2    0
1    251    0    1    0
1    254    0    1    0
1    63    0    2    0
1    25    0    2    0
1    197    0    1    0
1    206    0    1    0
1    100    0    2    0
1    124    0    2    0
1    43    0    2    0
1    54    0    2    0
1    127    0    2    0
1    15    0    2    0
1    661    0    2    0
1    196    0    1    0
1    2072    0    2    0
1    76    0    2    0
1    192    0    1    0
1    1971    0    2    0
1    2104    0    2    0
1    11    0    2    0
1    73    0    2    0
1    2678    0    2    0
1    269    0    1    0
1    135    0    2    0
1    2435    0    2    0
1    190    0    1    0
1    202    0    1    0
1    270    0    1    0
1    66    0    2    0
1    182    0    1    0
1    247    0    1    0
1    2430    0    2    0
1    241    0    1    0
1    79    0    2    0
1    177    0    1    0
1    61    0    2    0
1    53    0    2    0
1    60    0    2    0
1    5    0    2    0
1    47    0    2    0
1    72    0    2    0
1    2106    0    2    0
1    543    0    2    0
1    2066    0    2    0
1    199    0    1    0
1    215    0    1    0
1    255    0    1    0
1    28    0    2    0
1    119    0    2    0
1    262    0    1    0
1    276    0    1    0
1    99    0    2    0
1    129    0    2    0
1    253    0    1    0
1    115    0    2    0
1    55    0    2    0
1    116    0    2    0
1    212    0    1    0
1    2474    0    2    0
1    452    0    2    0
1    7    0    2    0
1    40    0    2    0
1    201    0    1    0
1    29    0    2    0
1    2096    0    2    0
1    114    0    2    0
1    179    0    1    0
1    132    0    2    0
1    186    0    1    0
1    198    0    1    0
1    244    0    1    0
1    69    0    2    0
1    193    0    1    0
1    93    0    2    0
1    249    0    1    0
1    209    0    1    0
1    92    0    2    0
1    272    0    1    0
1    2067    0    2    0
1    2084    0    2    0
1    2105    0    2    0
1    139    0    2    0
1    2    0    2    0
1    559    0    2    0
1    651    0    2    0
1    107    0    2    0
1    208    0    1    0
1    82    0    2    0
1    1976    0    2    0
1    4    0    2    0
1    120    0    2    0
1    106    0    2    0
1    204    0    1    0
1    178    0    1    0
1    19    0    2    0
1    14    0    2    0
1    130    0    2    0
1    89    0    2    0
1    239    0    1    0
1    277    0    1    0
1    32    0    2    0
1    36    0    2    0
1    242    0    1    0
1    1961    0    2    0
1    1996    0    2    0
1    2454    0    2    0
1    200    0    1    0
1    174    0    1    0
1    1986    0    2    0
1    37    0    2    0
1    189    0    1    0
1    111    0    2    0
1    194    0    1    0
1    185    0    1    0
1    250    0    1    0
1    1341    0    2    0
1    90    0    2    0
1    6    0    2    0
1    78    0    2    0
1    2078    0    2    0
1    211    0    1    0
1    210    0    1    0
1    275    0    1    0
1    49    0    2    0
1    65    0    2    0
1    169    0    1    0
1    252    0    1    0
1    123    0    2    0
3    350    1    0    1    452
3    335    1    0    1    452
3    409    1    0    1    452
0    546    7    1    2    1    3
0    560    5    1    1    559
3    369    1    0    1    1083
3    367    1    0    1    1083
0    1385    5    1    1    1384
3    411    1    0    1    2066
3    337    1    0    1    2066
3    384    1    0    1    2066
0    157    7    1    4    2090    2084    2078    2072
0    547    5    1    1    546
3    218    5    0    1    44
3    219    5    0    1    132
3    220    5    0    1    82
3    221    5    0    1    96
3    235    5    0    1    69
3    236    5    0    1    120
3    237    5    0    1    57
3    238    5    0    1    108
0    258    7    1    3    2    15    661
2    480    1    661
0    486    7    1    2    37    37
2    654    1    452
2    655    1    8
2    658    1    8
2    772    1    543
2    795    1    651
0    865    5    3    1    860
0    875    5    5    1    868
0    882    7    1    2    11    868
0    1251    7    2    4    132    82    96    44
0    1254    7    2    4    120    57    108    69
2    1261    1    543
2    1284    1    651
0    1344    5    3    1    1341
0    1351    5    3    1    1348
2    1394    1    2104
2    1418    1    2105
0    2433    5    1    1    2427
0    2434    5    1    1    2430
0    2441    5    1    1    2435
0    2442    5    1    1    2438
0    2449    5    1    1    2443
0    2450    5    1    1    2446
0    2478    5    1    1    2474
2    1631    1    2104
2    1655    1    2105
2    1710    1    16
2    1721    1    16
0    2682    5    1    1    2678
0    1955    7    3    2    7    661
0    1959    5    3    1    1956
0    1964    5    3    1    1961
0    1969    5    3    1    1966
0    1974    5    3    1    1971
0    1979    5    3    1    1976
0    1984    5    3    1    1981
0    1989    5    3    1    1986
0    1994    5    3    1    1991
0    1999    5    5    1    1996
2    2001    1    29
2    2012    1    29
0    2070    5    5    1    2067
0    2076    5    3    1    2072
0    2082    5    3    1    2078
0    2088    5    3    1    2084
0    2094    5    3    1    2090
0    2099    5    2    1    2096
0    2103    5    2    1    2100
0    2457    5    1    1    2451
0    2458    5    1    1    2454
2    2461    1    1348
2    2464    1    1341
2    2471    1    1956
2    2479    1    1966
2    2482    1    1961
2    2487    1    1976
2    2490    1    1971
2    2495    1    1986
2    2498    1    1981
2    2505    1    1996
2    2508    1    1991
2    2675    1    2067
2    2683    1    2078
2    2686    1    2072
2    2691    1    2090
2    2694    1    2084
2    2699    1    2100
2    2702    1    2096
3    158    5    0    1    157
3    259    5    0    1    258
0    487    5    2    1    486
3    391    1    0    1    654
0    1475    6    1    2    2430    2433
0    1476    6    1    2    2427    2434
0    1484    6    1    2    2438    2441
0    1485    6    1    2    2435    2442
0    1493    6    1    2    2446    2449
0    1494    6    1    2    2443    2450
0    2459    6    1    2    2454    2457
0    2460    6    1    2    2451    2458
3    173    7    0    2    94    654
0    216    7    1    2    2106    1955
3    223    5    0    1    1955
3    234    6    0    2    567    1955
0    1253    5    1    1    1251
0    1256    5    1    1    1254
0    558    7    2    2    1254    1251
2    748    1    655
0    784    5    10    1    772
0    807    5    10    1    795
0    821    7    1    3    80    772    795
0    825    7    1    3    68    772    795
0    829    7    1    3    79    772    795
0    833    7    1    3    78    772    795
0    837    7    1    3    77    772    795
0    881    7    1    2    11    875
2    994    1    655
0    1273    5    10    1    1261
0    1296    5    10    1    1284
0    1310    7    1    3    76    1261    1284
0    1314    7    1    3    75    1261    1284
0    1318    7    1    3    74    1261    1284
0    1322    7    1    3    73    1261    1284
0    1326    7    1    3    72    1261    1284
0    1406    5    10    1    1394
0    1430    5    10    1    1418
0    1444    7    1    3    114    1394    1418
0    1448    7    1    3    113    1394    1418
0    1452    7    1    3    112    1394    1418
0    1456    7    1    3    111    1394    1418
0    1460    7    1    2    1394    1418
0    1477    6    3    2    1475    1476
0    1486    6    3    2    1484    1485
0    1495    6    2    2    1493    1494
0    2477    5    1    1    2471
0    1499    6    1    2    2471    2478
0    2485    5    1    1    2479
0    2486    5    1    1    2482
0    2493    5    1    1    2487
0    2494    5    1    1    2490
0    1643    5    10    1    1631
0    1667    5    10    1    1655
0    1681    7    1    3    118    1631    1655
0    1685    7    1    3    107    1631    1655
0    1689    7    1    3    117    1631    1655
0    1693    7    1    3    116    1631    1655
0    1697    7    1    3    115    1631    1655
0    1716    5    4    1    1710
0    1728    5    5    1    1721
0    2681    5    1    1    2675
0    1776    6    1    2    2675    2682
0    2689    5    1    1    2683
0    2690    5    1    1    2686
0    2697    5    1    1    2691
0    2698    5    1    1    2694
2    1831    1    658
2    1893    1    658
0    2007    5    4    1    2001
0    2018    5    4    1    2012
0    2467    5    1    1    2461
0    2468    5    1    1    2464
0    2501    5    1    1    2495
0    2502    5    1    1    2498
0    2511    5    1    1    2505
0    2512    5    1    1    2508
0    2518    6    2    2    2459    2460
2    2551    1    1344
2    2559    1    1351
2    2567    1    1959
2    2575    1    1964
2    2583    1    1969
2    2591    1    1974
2    2599    1    1979
2    2607    1    1984
2    2615    1    1989
2    2623    1    1994
0    2705    5    1    1    2699
0    2706    5    1    1    2702
2    2735    1    1999
2    2743    1    2070
2    2751    1    2076
2    2759    1    2082
2    2767    1    2088
2    2775    1    2094
3    217    5    0    1    216
0    550    7    1    2    2106    1253
0    552    7    1    2    567    1256
3    325    1    0    1    558
0    894    3    1    2    881    882
0    1498    6    1    2    2474    2477
0    1507    6    1    2    2482    2485
0    1508    6    1    2    2479    2486
0    1516    6    1    2    2490    2493
0    1517    6    1    2    2487    2494
0    1775    6    1    2    2678    2681
0    1784    6    1    2    2686    2689
0    1785    6    1    2    2683    2690
0    1793    6    1    2    2694    2697
0    1794    6    1    2    2691    2698
0    2469    6    1    2    2464    2467
0    2470    6    1    2    2461    2468
0    2503    6    1    2    2498    2501
0    2504    6    1    2    2495    2502
0    2513    6    1    2    2508    2511
0    2514    6    1    2    2505    2512
0    2707    6    1    2    2702    2705
0    2708    6    1    2    2699    2706
3    261    5    0    1    558
0    551    5    1    1    550
0    553    5    1    1    552
0    818    7    1    3    93    784    807
0    819    7    1    3    55    772    807
0    820    7    1    3    67    784    795
0    822    7    1    3    81    784    807
0    823    7    1    3    43    772    807
0    824    7    1    3    56    784    795
0    826    7    1    3    92    784    807
0    827    7    1    3    54    772    807
0    828    7    1    3    66    784    795
0    830    7    1    3    91    784    807
0    831    7    1    3    53    772    807
0    832    7    1    3    65    784    795
0    834    7    1    3    90    784    807
0    835    7    1    3    52    772    807
0    836    7    1    3    64    784    795
0    1307    7    1    3    89    1273    1296
0    1308    7    1    3    51    1261    1296
0    1309    7    1    3    63    1273    1284
0    1311    7    1    3    88    1273    1296
0    1312    7    1    3    50    1261    1296
0    1313    7    1    3    62    1273    1284
0    1315    7    1    3    87    1273    1296
0    1316    7    1    3    49    1261    1296
0    1317    7    1    2    1273    1284
0    1319    7    1    3    86    1273    1296
0    1320    7    1    3    48    1261    1296
0    1321    7    1    3    61    1273    1284
0    1323    7    1    3    85    1273    1296
0    1324    7    1    3    47    1261    1296
0    1325    7    1    3    60    1273    1284
0    1441    7    1    3    138    1406    1430
0    1442    7    1    3    102    1394    1430
0    1443    7    1    3    126    1406    1418
0    1445    7    1    3    137    1406    1430
0    1446    7    1    3    101    1394    1430
0    1447    7    1    3    125    1406    1418
0    1449    7    1    3    136    1406    1430
0    1450    7    1    3    100    1394    1430
0    1451    7    1    3    124    1406    1418
0    1453    7    1    3    135    1406    1430
0    1454    7    1    3    99    1394    1430
0    1455    7    1    3    123    1406    1418
0    1457    7    1    2    1406    1430
0    1458    7    1    2    1394    1430
0    1459    7    1    2    1406    1418
0    1481    5    2    1    1477
0    1490    5    2    1    1486
0    1500    6    3    2    1498    1499
0    1509    6    3    2    1507    1508
0    1518    6    2    2    1516    1517
2    1521    1    1495
2    1525    1    1495
0    2557    5    1    1    2551
0    2565    5    1    1    2559
0    2573    5    1    1    2567
0    2581    5    1    1    2575
0    2589    5    1    1    2583
0    2597    5    1    1    2591
0    2605    5    1    1    2599
0    2613    5    1    1    2607
0    2621    5    1    1    2615
0    2629    5    1    1    2623
0    1678    7    1    3    142    1643    1667
0    1679    7    1    3    106    1631    1667
0    1680    7    1    3    130    1643    1655
0    1682    7    1    3    131    1643    1667
0    1683    7    1    3    95    1631    1667
0    1684    7    1    3    119    1643    1655
0    1686    7    1    3    141    1643    1667
0    1687    7    1    3    105    1631    1667
0    1688    7    1    3    129    1643    1655
0    1690    7    1    3    140    1643    1667
0    1691    7    1    3    104    1631    1667
0    1692    7    1    3    128    1643    1655
0    1694    7    1    3    139    1643    1667
0    1695    7    1    3    103    1631    1667
0    1696    7    1    3    127    1643    1655
0    1734    7    1    2    19    1716
0    1736    7    1    2    4    1716
0    1738    7    1    2    20    1716
0    1740    7    1    2    5    1716
0    1742    7    1    2    21    1728
0    1744    7    1    2    22    1728
0    1746    7    1    2    23    1728
0    1748    7    1    2    6    1728
0    1750    7    1    2    24    1728
0    1777    6    3    2    1775    1776
0    1786    6    3    2    1784    1785
0    1795    6    2    2    1793    1794
0    2023    7    1    2    25    2007
0    2025    7    1    2    32    2007
0    2027    7    1    2    26    2007
0    2029    7    1    2    33    2007
0    2031    7    1    2    27    2018
0    2033    7    1    2    34    2018
0    2035    7    1    2    35    2018
0    2037    7    1    2    28    2018
0    2741    5    1    1    2735
0    2749    5    1    1    2743
0    2757    5    1    1    2751
0    2765    5    1    1    2759
0    2773    5    1    1    2767
0    2781    5    1    1    2775
0    2515    6    2    2    2469    2470
0    2522    5    1    1    2518
0    2525    6    2    2    2513    2514
0    2528    6    2    2    2503    2504
0    2730    6    2    2    2707    2708
0    554    7    4    2    551    553
0    838    3    3    4    818    819    820    821
0    841    3    5    4    822    823    824    825
0    846    3    5    4    826    827    828    829
0    854    3    2    4    830    831    832    833
0    857    3    3    4    834    835    836    837
0    1327    3    4    4    1307    1308    1309    1310
0    1329    3    3    4    1311    1312    1313    1314
0    1331    3    2    4    1315    1316    1317    1318
0    1333    3    2    4    1319    1320    1321    1322
0    1335    3    2    4    1323    1324    1325    1326
0    1461    3    4    4    1441    1442    1443    1444
0    1464    3    4    4    1445    1446    1447    1448
0    1467    3    3    4    1449    1450    1451    1452
0    1470    3    4    4    1453    1454    1455    1456
0    1473    3    3    4    1457    1458    1459    1460
0    1698    3    4    4    1682    1683    1684    1685
0    1701    3    4    4    1686    1687    1688    1689
0    1704    3    3    4    1690    1691    1692    1693
0    1707    3    2    4    1694    1695    1696    1697
0    2634    3    2    4    1678    1679    1680    1681
3    319    1    0    1    554
0    1504    5    2    1    1500
0    1513    5    2    1    1509
0    1524    5    1    1    1521
0    1528    5    1    1    1525
2    1529    1    1518
2    1533    1    1518
0    1538    7    1    3    1486    1477    1521
0    1541    7    1    3    1490    1481    1525
0    1781    5    2    1    1777
0    1790    5    2    1    1786
2    1806    1    1795
2    1810    1    1795
0    2734    5    1    1    2730
0    2521    5    1    1    2515
0    2524    6    1    2    2515    2522
0    2531    5    1    1    2525
0    2532    5    1    1    2528
0    144    7    1    2    838    860
0    147    7    1    2    846    860
0    152    7    1    2    841    860
3    160    5    0    1    1464
3    162    5    0    1    1467
3    164    5    0    1    1461
3    166    5    0    1    1329
3    168    5    0    1    1327
3    171    5    0    1    857
0    175    7    1    4    480    483    36    554
0    187    7    1    4    480    483    554    547
2    516    1    838
0    852    5    2    1    846
0    885    7    1    2    841    875
0    887    7    1    2    846    875
0    893    7    1    2    1327    868
0    1028    5    2    1    838
0    1031    5    4    1    841
0    1035    5    6    1    846
2    1041    1    854
2    1049    1    857
2    1057    1    1327
2    1060    1    1329
2    1066    1    1331
2    1072    1    1333
2    1078    1    1335
0    1213    6    2    2    2099    1470
0    1218    6    2    2    2103    1473
2    1250    1    1704
0    1387    7    2    2    1461    1385
0    1389    5    2    1    1464
0    1537    7    1    3    1481    1486    1524
0    1540    7    1    3    1477    1490    1528
0    1735    7    1    2    841    1710
0    1737    7    1    2    846    1710
0    1739    7    1    2    854    1710
0    1741    7    1    2    857    1710
0    1743    7    1    2    1327    1721
0    1745    7    1    2    1329    1721
0    1747    7    1    2    1331    1721
0    1749    7    1    2    1333    1721
0    1751    7    1    2    1335    1721
0    2638    5    1    1    2634
0    2024    7    1    2    1698    2001
0    2026    7    1    2    1701    2001
0    2028    7    1    2    1704    2001
0    2030    7    1    2    1707    2001
0    2032    7    1    2    1461    2012
0    2034    7    1    2    1464    2012
0    2036    7    1    2    1467    2012
0    2038    7    1    2    1470    2012
2    2154    1    841
0    2523    6    1    2    2518    2521
0    2533    6    1    2    2528    2531
0    2534    6    1    2    2525    2532
2    2631    1    1698
2    2639    1    1704
2    2642    1    1701
2    2647    1    1461
2    2650    1    1707
2    2655    1    1467
2    2658    1    1464
2    2665    1    1473
2    2668    1    1470
3    153    3    0    2    865    152
3    176    5    0    1    175
3    188    5    0    1    187
3    299    1    0    1    1041
3    301    1    0    1    1049
3    286    1    0    1    1057
3    303    1    0    1    1060
3    288    1    0    1    1066
3    305    1    0    1    1072
3    290    1    0    1    1078
0    1532    5    1    1    1529
0    1536    5    1    1    1533
0    1539    4    1    2    1537    1538
0    1542    4    1    2    1540    1541
0    1544    7    1    3    1509    1500    1529
0    1547    7    1    3    1513    1504    1533
0    2065    3    1    2    2037    2038
0    1809    5    1    1    1806
0    1813    5    1    1    1810
0    1821    7    1    3    1786    1777    1806
0    1824    7    1    3    1790    1781    1810
0    2538    6    2    2    2523    2524
0    2546    6    2    2    2533    2534
0    2554    3    2    2    1734    1735
0    2562    3    2    2    1736    1737
0    2570    3    2    2    1738    1739
0    2578    3    2    2    1740    1741
0    2586    3    2    2    1742    1743
0    2594    3    2    2    1744    1745
0    2602    3    2    2    1746    1747
0    2610    3    2    2    1748    1749
0    2618    3    2    2    1750    1751
0    2626    3    2    2    2023    2024
0    2738    3    2    2    2025    2026
0    2746    3    2    2    2027    2028
0    2754    3    2    2    2029    2030
0    2762    3    2    2    2031    2032
0    2770    3    2    2    2033    2034
0    2778    3    2    2    2035    2036
0    456    7    5    3    1389    1387    40
0    466    5    1    1    1387
0    562    6    4    2    560    852
0    883    7    1    2    516    875
0    889    7    1    2    1049    868
0    891    7    1    2    1041    875
0    1043    5    6    1    1041
0    1051    5    5    1    1049
0    1062    5    2    1    1060
0    1068    5    2    1    1066
0    1074    5    2    1    1072
0    1080    5    2    1    1078
0    1225    7    1    2    2099    1213
0    1227    7    1    2    1213    1470
0    1232    7    1    2    2103    1218
0    1234    7    1    2    1218    1473
0    1543    7    1    3    1504    1509    1532
0    1546    7    1    3    1500    1513    1536
0    2637    5    1    1    2631
0    1753    6    1    2    2631    2638
0    2645    5    1    1    2639
0    2646    5    1    1    2642
0    2653    5    1    1    2647
0    2654    5    1    1    2650
0    1820    7    1    3    1781    1786    1809
0    1823    7    1    3    1777    1790    1813
2    2107    1    1031
2    2110    1    1028
2    2118    1    1035
0    2123    5    2    1    1057
0    2151    5    2    1    852
0    2158    5    1    1    2154
2    2161    1    1031
2    2164    1    1028
2    2172    1    1035
2    2235    1    516
2    2262    1    1035
2    2350    1    1035
0    2535    6    2    2    1542    1539
0    2661    5    1    1    2655
0    2662    5    1    1    2658
0    2671    5    1    1    2665
0    2672    5    1    1    2668
0    468    7    2    3    40    1389    466
0    897    3    2    2    887    889
0    898    3    2    2    891    893
0    1228    3    2    2    1225    1227
0    1235    3    2    2    1232    1234
0    1545    4    1    2    1543    1544
0    1548    4    1    2    1546    1547
0    2542    5    1    1    2538
0    2550    5    1    1    2546
0    1561    6    1    2    2554    2557
0    2558    5    1    1    2554
0    1565    6    1    2    2562    2565
0    2566    5    1    1    2562
0    1569    6    1    2    2570    2573
0    2574    5    1    1    2570
0    1573    6    1    2    2578    2581
0    2582    5    1    1    2578
0    1577    6    1    2    2586    2589
0    2590    5    1    1    2586
0    1581    6    1    2    2594    2597
0    2598    5    1    1    2594
0    1585    6    1    2    2602    2605
0    2606    5    1    1    2602
0    1589    6    1    2    2610    2613
0    2614    5    1    1    2610
0    1593    6    1    2    2618    2621
0    2622    5    1    1    2618
0    1597    6    1    2    2626    2629
0    2630    5    1    1    2626
0    1752    6    1    2    2634    2637
0    1761    6    1    2    2642    2645
0    1762    6    1    2    2639    2646
0    1770    6    1    2    2650    2653
0    1771    6    1    2    2647    2654
0    1822    4    1    2    1820    1821
0    1825    4    1    2    1823    1824
0    2039    6    1    2    2738    2741
0    2742    5    1    1    2738
0    2043    6    1    2    2746    2749
0    2750    5    1    1    2746
0    2047    6    1    2    2754    2757
0    2758    5    1    1    2754
0    2051    6    1    2    2762    2765
0    2766    5    1    1    2762
0    2055    6    1    2    2770    2773
0    2774    5    1    1    2770
0    2059    6    1    2    2778    2781
0    2782    5    1    1    2778
0    2663    6    1    2    2658    2661
0    2664    6    1    2    2655    2662
0    2673    6    1    2    2668    2671
0    2674    6    1    2    2665    2672
0    146    7    1    2    562    865
0    462    5    2    1    456
0    2113    5    1    1    2107
0    2114    5    1    1    2110
0    2122    5    1    1    2118
0    2129    5    1    1    2123
2    592    1    562
0    2167    5    1    1    2161
0    2168    5    1    1    2164
0    2176    5    1    1    2172
0    2241    5    1    1    2235
0    2266    5    1    1    2262
0    743    5    4    1    456
2    749    1    456
0    886    7    1    2    562    868
3    284    1    0    1    897
3    321    1    0    1    897
3    297    1    0    1    898
3    280    1    0    1    898
2    995    1    456
0    1006    5    4    1    456
0    1550    6    1    2    2535    2542
0    2354    5    1    1    2350
0    2541    5    1    1    2535
0    1562    6    1    2    2551    2558
0    1566    6    1    2    2559    2566
0    1570    6    1    2    2567    2574
0    1574    6    1    2    2575    2582
0    1578    6    1    2    2583    2590
0    1582    6    1    2    2591    2598
0    1586    6    1    2    2599    2606
0    1590    6    1    2    2607    2614
0    1594    6    1    2    2615    2622
0    1598    6    1    2    2623    2630
0    1754    6    3    2    1752    1753
0    1763    6    3    2    1761    1762
0    1772    6    2    2    1770    1771
0    2040    6    1    2    2735    2742
0    2044    6    1    2    2743    2750
0    2048    6    1    2    2751    2758
0    2052    6    1    2    2759    2766
0    2056    6    1    2    2767    2774
0    2060    6    1    2    2775    2782
2    2115    1    1043
2    2126    1    1051
2    2131    1    1068
2    2134    1    1062
2    2141    1    1080
2    2144    1    1074
0    2157    5    1    1    2151
0    2160    6    1    2    2151    2158
2    2169    1    1043
2    2177    1    1068
2    2180    1    1062
2    2187    1    1080
2    2190    1    1074
0    2207    5    2    1    562
2    2254    1    1043
2    2334    1    1051
2    2342    1    1043
2    2422    1    1051
0    2543    6    2    2    1548    1545
0    2709    6    2    2    2673    2674
0    2712    6    2    2    2663    2664
0    2727    6    2    2    1825    1822
3    148    3    0    2    146    147
0    569    6    1    2    2110    2113
0    570    6    1    2    2107    2114
0    599    6    1    2    2164    2167
0    600    6    1    2    2161    2168
0    896    3    2    2    885    886
0    1549    6    1    2    2538    2541
0    1243    5    2    1    1228
0    1245    5    2    1    1235
2    1257    1    468
2    1258    1    468
0    1563    6    1    2    1561    1562
0    1567    6    1    2    1565    1566
0    1571    6    1    2    1569    1570
0    1575    6    1    2    1573    1574
0    1579    6    1    2    1577    1578
0    1583    6    1    2    1581    1582
0    1587    6    1    2    1585    1586
0    1591    6    1    2    1589    1590
0    1595    6    1    2    1593    1594
0    1599    6    1    2    1597    1598
0    2041    6    1    2    2039    2040
0    2045    6    1    2    2043    2044
0    2049    6    1    2    2047    2048
0    2053    6    1    2    2051    2052
0    2057    6    1    2    2055    2056
0    2061    6    1    2    2059    2060
0    2159    6    1    2    2154    2157
2    475    1    462
0    490    7    1    2    1078    743
0    496    7    1    2    1698    743
0    502    7    1    2    1701    743
0    508    7    1    2    1250    743
0    765    7    1    2    1057    749
0    769    7    1    2    1060    749
0    571    6    3    2    569    570
0    2121    5    1    1    2115
0    579    6    1    2    2115    2122
0    587    6    1    2    2126    2129
0    2130    5    1    1    2126
0    596    5    2    1    592
0    601    6    3    2    599    600
0    2175    5    1    1    2169
0    609    6    1    2    2169    2176
0    2258    5    1    1    2254
0    1014    7    1    2    1057    995
0    1018    7    1    2    1060    995
0    717    7    1    2    1078    1006
0    723    7    1    2    1698    1006
0    729    7    1    2    1701    1006
0    735    7    1    2    1250    1006
0    753    5    4    1    749
3    282    1    0    1    896
3    323    1    0    1    896
0    2338    5    1    1    2334
0    999    5    4    1    995
0    1091    6    1    2    1549    1550
0    2346    5    1    1    2342
0    2426    5    1    1    2422
2    1337    1    462
0    2549    5    1    1    2543
0    1552    6    1    2    2543    2550
0    1600    5    1    1    1599
0    1596    5    1    1    1595
0    1592    5    1    1    1591
0    1588    5    1    1    1587
0    1584    5    1    1    1583
0    1580    5    1    1    1579
0    1576    5    1    1    1575
0    1572    5    1    1    1571
0    1568    5    1    1    1567
0    1564    5    1    1    1563
0    2062    5    1    1    2061
0    2058    5    1    1    2057
0    2054    5    1    1    2053
0    2050    5    1    1    2049
0    2046    5    1    1    2045
0    2042    5    1    1    2041
0    1758    5    2    1    1754
0    1767    5    2    1    1763
2    1798    1    1772
2    1802    1    1772
0    2733    5    1    1    2727
0    1829    6    1    2    2727    2734
0    2137    5    1    1    2131
0    2138    5    1    1    2134
0    2147    5    1    1    2141
0    2148    5    1    1    2144
0    2183    5    1    1    2177
0    2184    5    1    1    2180
0    2193    5    1    1    2187
0    2194    5    1    1    2190
0    2210    6    2    2    2159    2160
0    2213    5    1    1    2207
0    2715    5    1    1    2709
0    2716    5    1    1    2712
0    1094    7    1    2    1235    1245
0    1096    7    1    2    1228    1243
0    578    6    1    2    2118    2121
0    588    6    1    2    2123    2130
0    608    6    1    2    2172    2175
2    742    1    1257
2    1005    1    1257
0    1092    5    1    1    1091
0    1551    6    1    2    2546    2549
0    1554    7    1    5    1600    1596    1592    1588    1584
0    1555    7    1    5    1580    1576    1572    1568    1564
0    1557    7    1    2    2065    2062
0    1558    7    1    5    2058    2054    2050    2046    2042
0    1828    6    1    2    2730    2733
2    1845    1    1258
2    1907    1    1258
0    2139    6    1    2    2134    2137
0    2140    6    1    2    2131    2138
0    2149    6    1    2    2144    2147
0    2150    6    1    2    2141    2148
0    2185    6    1    2    2180    2183
0    2186    6    1    2    2177    2184
0    2195    6    1    2    2190    2193
0    2196    6    1    2    2187    2194
0    2717    6    1    2    2712    2715
0    2718    6    1    2    2709    2716
0    154    3    1    2    1094    1245
0    155    3    1    2    1096    1243
0    763    7    1    2    1057    753
0    767    7    1    2    1060    753
0    531    7    1    2    1066    753
0    537    7    1    2    1072    753
0    575    5    2    1    571
0    580    6    3    2    578    579
0    589    6    2    2    587    588
0    605    5    2    1    601
0    610    6    2    2    608    609
0    1012    7    1    2    1057    999
0    1016    7    1    2    1060    999
0    705    7    1    2    1066    999
0    711    7    1    2    1072    999
0    1093    7    2    2    1092    14
2    1355    1    475
0    1553    6    2    2    1551    1552
0    1556    7    1    2    1554    1555
0    1559    7    1    2    1557    1558
2    1601    1    1337
0    1801    5    1    1    1798
0    1805    5    1    1    1802
0    1815    7    1    3    1763    1754    1798
0    1818    7    1    3    1767    1758    1802
0    1830    6    2    2    1828    1829
2    1836    1    475
2    1850    1    475
2    1898    1    1337
2    1912    1    1337
0    2197    6    2    2    2149    2150
0    2200    6    2    2    2139    2140
0    2214    5    1    1    2210
0    2215    6    1    2    2210    2213
0    2217    6    2    2    2195    2196
0    2220    6    2    2    2185    2186
0    2722    6    2    2    2717    2718
3    156    6    0    2    154    155
0    492    7    1    2    490    742
0    498    7    1    2    496    742
0    504    7    1    2    502    742
0    510    7    1    2    508    742
0    519    3    1    2    763    765
0    525    3    1    2    767    769
0    533    7    1    2    531    748
0    539    7    1    2    537    748
0    693    3    1    2    1012    1014
0    699    3    1    2    1016    1018
0    707    7    1    2    705    994
0    713    7    1    2    711    994
0    719    7    1    2    717    1005
0    725    7    1    2    723    1005
0    731    7    1    2    729    1005
0    737    7    1    2    735    1005
3    401    1    0    1    1093
0    1560    7    2    3    1556    1559    894
0    1814    7    1    3    1758    1763    1801
0    1817    7    1    3    1754    1767    1805
0    2216    6    1    2    2207    2214
3    227    5    0    1    1830
3    229    5    0    1    1553
0    493    5    2    1    492
0    499    5    2    1    498
0    505    5    2    1    504
0    511    5    2    1    510
0    521    7    1    2    519    748
0    527    7    1    2    525    748
0    534    5    2    1    533
0    540    5    2    1    539
0    584    5    2    1    580
2    613    1    589
2    617    1    589
2    621    1    610
2    625    1    610
0    676    7    1    2    1344    1355
0    695    7    1    2    693    994
0    701    7    1    2    699    994
0    708    5    2    1    707
0    714    5    2    1    713
0    720    5    2    1    719
0    726    5    2    1    725
0    732    5    2    1    731
0    738    5    2    1    737
0    1087    5    1    1    1093
0    1108    7    1    2    1344    1601
0    1361    5    4    1    1355
0    1369    7    1    2    1351    1355
0    1373    7    1    2    1959    1355
0    1377    7    1    2    1964    1355
3    311    1    0    1    1560
0    1607    5    4    1    1601
0    1615    7    1    2    1351    1601
0    1619    7    1    2    1959    1601
0    1623    7    1    2    1964    1601
0    1816    4    1    2    1814    1815
0    1819    4    1    2    1817    1818
0    2726    5    1    1    2722
0    1842    5    2    1    1836
0    1858    7    1    2    1969    1836
0    1863    7    1    2    1974    1836
0    1866    7    1    2    1979    1836
0    1868    7    1    2    1984    1836
0    1870    7    1    2    1989    1850
0    1872    7    1    2    1994    1850
0    1874    7    1    2    1999    1850
0    1876    7    1    2    2070    1850
0    1904    5    2    1    1898
0    1920    7    1    2    1969    1898
0    1925    7    1    2    1974    1898
0    1928    7    1    2    1979    1898
0    1930    7    1    2    1984    1898
0    1932    7    1    2    1989    1912
0    1934    7    1    2    1994    1912
0    1936    7    1    2    1999    1912
0    1938    7    1    2    2070    1912
0    2203    5    1    1    2197
0    2204    5    1    1    2200
0    2223    5    1    1    2217
0    2224    5    1    1    2220
0    2238    6    2    2    2215    2216
3    150    5    0    1    1560
0    522    5    2    1    521
0    528    5    2    1    527
0    696    5    2    1    695
0    702    5    2    1    701
0    1881    7    2    2    1866    1831
0    1883    7    2    2    1868    1831
0    1885    7    2    2    1870    1845
0    1887    7    2    2    1872    1845
0    1889    7    2    2    1874    1845
0    1891    7    2    2    1876    1845
0    1943    7    2    2    1928    1893
0    1945    7    2    2    1930    1893
0    1947    7    2    2    1932    1907
0    1949    7    2    2    1934    1907
0    1951    7    2    2    1936    1907
0    1953    7    2    2    1938    1907
0    2205    6    1    2    2200    2203
0    2206    6    1    2    2197    2204
0    2225    6    1    2    2220    2223
0    2226    6    1    2    2217    2224
0    2719    6    2    2    1819    1816
0    616    5    1    1    613
0    620    5    1    1    617
0    624    5    1    1    621
0    628    5    1    1    625
0    630    7    1    3    580    571    613
0    633    7    1    3    584    575    617
0    636    7    1    3    601    592    621
0    639    7    1    3    605    596    625
0    645    6    1    2    2238    2241
0    2242    5    1    1    2238
0    675    7    1    2    1999    1361
0    1107    7    1    2    1999    1607
0    1368    7    1    2    2070    1361
0    1371    7    1    2    2076    1361
0    1375    7    1    2    2082    1361
0    1614    7    1    2    2070    1607
0    1617    7    1    2    2076    1607
0    1621    7    1    2    2082    1607
0    1856    7    1    2    2088    1842
0    1861    7    1    2    2094    1842
0    1918    7    1    2    2088    1904
0    1923    7    1    2    2094    1904
0    2230    6    2    2    2205    2206
0    2246    6    2    2    2225    2226
2    2270    1    511
2    2278    1    505
2    2286    1    499
2    2294    1    493
2    2302    1    540
2    2310    1    534
2    2358    1    738
2    2366    1    732
2    2374    1    726
2    2382    1    720
2    2390    1    714
2    2398    1    708
0    629    7    1    3    575    580    616
0    632    7    1    3    571    584    620
0    635    7    1    3    596    601    624
0    638    7    1    3    592    605    628
0    646    6    1    2    2235    2242
0    677    3    1    2    675    676
0    1827    6    1    2    2719    2726
0    907    7    1    2    1891    511
0    915    7    1    2    1889    505
0    922    7    1    2    1887    499
0    924    7    1    2    493    1885
0    937    7    1    2    1883    540
0    946    7    1    2    1881    534
0    1109    3    1    2    1107    1108
0    1125    7    1    2    1953    738
0    1133    7    1    2    1951    732
0    1140    7    1    2    1949    726
0    1142    7    1    2    720    1947
0    1155    7    1    2    1945    714
0    1164    7    1    2    1943    708
0    1378    3    2    2    1368    1369
0    1380    3    2    2    1371    1373
0    1382    3    2    2    1375    1377
0    1624    3    2    2    1614    1615
0    1626    3    2    2    1617    1619
0    1628    3    2    2    1621    1623
0    2725    5    1    1    2719
0    1859    3    1    2    1856    1858
0    1864    3    1    2    1861    1863
0    1921    3    1    2    1918    1920
0    1926    3    1    2    1923    1925
2    2267    1    1891
2    2275    1    1889
2    2283    1    1887
2    2291    1    1885
2    2299    1    1883
2    2307    1    1881
2    2318    1    528
2    2326    1    522
2    2355    1    1953
2    2363    1    1951
2    2371    1    1949
2    2379    1    1947
2    2387    1    1945
2    2395    1    1943
2    2406    1    702
2    2414    1    696
0    647    6    1    2    645    646
0    631    4    1    2    629    630
0    634    4    1    2    632    633
0    637    4    1    2    635    636
0    640    4    1    2    638    639
0    2234    5    1    1    2230
0    2250    5    1    1    2246
0    679    7    1    2    677    1031
0    1826    6    1    2    2722    2725
0    2274    5    1    1    2270
0    2282    5    1    1    2278
0    2290    5    1    1    2286
0    2298    5    1    1    2294
0    2306    5    1    1    2302
0    2314    5    1    1    2310
0    1110    7    1    2    1109    1031
0    2362    5    1    1    2358
0    2370    5    1    1    2366
0    2378    5    1    1    2374
0    2386    5    1    1    2382
0    2394    5    1    1    2390
0    2402    5    1    1    2398
0    1877    7    2    2    1859    1831
0    1879    7    2    2    1864    1831
0    1939    7    2    2    1921    1893
0    1941    7    2    2    1926    1893
0    143    7    1    2    647    865
0    671    7    1    2    1380    1043
0    674    7    1    2    1378    1035
0    686    6    1    2    1826    1827
0    2273    5    1    1    2267
0    900    6    1    2    2267    2274
0    2281    5    1    1    2275
0    909    6    1    2    2275    2282
0    2289    5    1    1    2283
0    917    6    1    2    2283    2290
0    2297    5    1    1    2291
0    926    6    1    2    2291    2298
0    2305    5    1    1    2299
0    929    6    1    2    2299    2306
0    2313    5    1    1    2307
0    939    6    1    2    2307    2314
0    2322    5    1    1    2318
0    2330    5    1    1    2326
0    967    7    1    2    1382    1051
0    1104    7    1    2    1626    1043
0    1106    7    1    2    1624    1035
0    2361    5    1    1    2355
0    1118    6    1    2    2355    2362
0    2369    5    1    1    2363
0    1127    6    1    2    2363    2370
0    2377    5    1    1    2371
0    1135    6    1    2    2371    2378
0    2385    5    1    1    2379
0    1144    6    1    2    2379    2386
0    2393    5    1    1    2387
0    1147    6    1    2    2387    2394
0    2401    5    1    1    2395
0    1157    6    1    2    2395    2402
0    2410    5    1    1    2406
0    2418    5    1    1    2414
0    1184    7    1    2    1628    1051
0    2227    6    2    2    634    631
0    2243    6    2    2    640    637
2    2251    1    1380
2    2259    1    1378
2    2331    1    1382
2    2339    1    1626
2    2347    1    1624
2    2419    1    1628
3    145    3    0    2    143    144
0    687    5    1    1    686
0    899    6    1    2    2270    2273
0    908    6    1    2    2278    2281
0    916    6    1    2    2286    2289
0    925    6    1    2    2294    2297
0    928    6    1    2    2302    2305
0    938    6    1    2    2310    2313
0    954    7    1    2    1879    528
0    961    7    1    2    1877    522
0    1117    6    1    2    2358    2361
0    1126    6    1    2    2366    2369
0    1134    6    1    2    2374    2377
0    1143    6    1    2    2382    2385
0    1146    6    1    2    2390    2393
0    1156    6    1    2    2398    2401
0    1172    7    1    2    1941    702
0    1179    7    1    2    1939    696
2    2315    1    1879
2    2323    1    1877
2    2403    1    1941
2    2411    1    1939
0    2233    5    1    1    2227
0    642    6    1    2    2227    2234
0    2249    5    1    1    2243
0    649    6    1    2    2243    2250
0    2257    5    1    1    2251
0    665    6    1    2    2251    2258
0    684    6    1    2    2259    2266
0    2265    5    1    1    2259
0    688    7    2    2    687    487
0    901    6    4    2    899    900
0    910    6    3    2    908    909
0    918    6    2    2    916    917
0    927    6    1    2    925    926
0    930    6    5    2    928    929
0    940    6    4    2    938    939
0    2337    5    1    1    2331
0    963    6    1    2    2331    2338
0    2345    5    1    1    2339
0    1099    6    1    2    2339    2346
0    1115    6    1    2    2347    2354
0    2353    5    1    1    2347
0    1119    6    4    2    1117    1118
0    1128    6    3    2    1126    1127
0    1136    6    2    2    1134    1135
0    1145    6    1    2    1143    1144
0    1148    6    5    2    1146    1147
0    1158    6    4    2    1156    1157
0    2425    5    1    1    2419
0    1181    6    1    2    2419    2426
0    641    6    1    2    2230    2233
0    648    6    1    2    2246    2249
0    664    6    1    2    2254    2257
0    683    6    1    2    2262    2265
3    395    1    0    1    688
0    2321    5    1    1    2315
0    948    6    1    2    2315    2322
0    2329    5    1    1    2323
0    956    6    1    2    2323    2330
0    962    6    1    2    2334    2337
0    1098    6    1    2    2342    2345
0    1114    6    1    2    2350    2353
0    2409    5    1    1    2403
0    1166    6    1    2    2403    2410
0    2417    5    1    1    2411
0    1174    6    1    2    2411    2418
0    1180    6    1    2    2422    2425
0    643    6    1    2    641    642
0    650    6    1    2    648    649
0    666    6    2    2    664    665
0    681    6    1    2    683    684
0    690    5    1    1    688
0    947    6    1    2    2318    2321
0    955    6    1    2    2326    2329
0    964    6    1    2    962    963
0    968    7    1    4    910    927    918    901
0    970    7    1    2    901    915
0    971    7    1    3    910    901    922
0    972    7    1    4    918    901    924    910
0    978    7    1    2    930    946
0    979    7    1    3    940    930    954
0    1100    6    2    2    1098    1099
0    1112    6    1    2    1114    1115
0    1165    6    1    2    2406    2409
0    1173    6    1    2    2414    2417
0    1182    6    1    2    1180    1181
0    1185    7    1    4    1128    1145    1136    1119
0    1187    7    1    2    1119    1133
0    1188    7    1    3    1128    1119    1140
0    1189    7    1    4    1136    1119    1142    1128
0    1195    7    1    2    1148    1164
0    1196    7    1    3    1158    1148    1172
0    644    5    1    1    643
0    884    7    1    2    650    868
0    949    6    3    2    947    948
0    957    6    2    2    955    956
0    969    5    1    1    968
0    973    3    2    4    907    970    971    972
0    1167    6    3    2    1165    1166
0    1175    6    2    2    1173    1174
0    1186    5    1    1    1185
0    1190    3    2    4    1125    1187    1188    1189
0    680    7    1    2    666    674
0    682    7    1    3    681    666    679
0    895    3    2    2    883    884
0    1025    7    2    2    644    487
0    1111    7    1    2    1100    1106
0    1113    7    1    3    1112    1100    1110
0    685    3    1    3    671    680    682
3    295    1    0    1    895
3    331    1    0    1    895
0    976    5    1    1    973
0    977    7    1    5    940    964    949    930    957
0    980    7    1    4    949    930    961    940
0    981    7    1    5    957    949    930    967    940
3    397    1    0    1    1025
0    1116    3    1    3    1104    1111    1113
0    1193    5    1    1    1190
0    1194    7    1    5    1158    1182    1167    1148    1175
0    1197    7    1    4    1167    1148    1179    1158
0    1198    7    1    5    1175    1167    1148    1184    1158
0    982    3    1    5    937    978    979    980    981
0    983    7    1    2    977    685
0    988    6    1    2    976    969
0    1027    5    1    1    1025
0    1199    3    1    5    1155    1195    1196    1197    1198
0    1200    7    1    2    1194    1116
0    1205    6    1    2    1193    1186
0    984    3    2    2    982    983
0    1085    7    1    3    690    1027    1830
0    1201    3    2    2    1199    1200
0    987    5    1    1    984
0    990    7    1    2    988    984
0    1204    5    1    1    1201
0    1207    7    1    2    1205    1201
0    989    7    1    2    973    987
0    1206    7    1    2    1190    1204
0    991    3    2    2    989    990
0    1208    3    3    2    1206    1207
3    329    1    0    1    1208
0    1221    6    2    2    1208    991
0    1238    7    1    2    1208    1221
0    1239    7    1    2    1221    991
0    1240    3    2    2    1238    1239
0    1247    5    2    1    1240
0    471    7    1    2    1240    1247
0    473    3    2    2    471    1247
3    231    5    0    1    473
0    1088    7    1    3    1553    1087    473
0    1089    7    2    3    1085    1088    554
3    308    1    0    1    1089
3    225    5    0    1    1089
3    274    0    0    0
3    266    0    0    0
3    191    0    0    0
3    265    0    0    0
3    268    0    0    0
3    264    0    0    0
3    271    0    0    0
3    184    0    0    0
3    213    0    0    0
3    273    0    0    0
3    214    0    0    0
3    203    0    0    0
3    181    0    0    0
3    240    0    0    0
3    207    0    0    0
3    205    0    0    0
3    267    0    0    0
3    278    0    0    0
3    256    0    0    0
3    246    0    0    0
3    257    0    0    0
3    183    0    0    0
3    279    0    0    0
3    180    0    0    0
3    263    0    0    0
3    195    0    0    0
3    245    0    0    0
3    243    0    0    0
3    248    0    0    0
3    251    0    0    0
3    254    0    0    0
3    197    0    0    0
3    206    0    0    0
3    196    0    0    0
3    192    0    0    0
3    269    0    0    0
3    190    0    0    0
3    202    0    0    0
3    270    0    0    0
3    182    0    0    0
3    247    0    0    0
3    241    0    0    0
3    177    0    0    0
3    199    0    0    0
3    215    0    0    0
3    255    0    0    0
3    262    0    0    0
3    276    0    0    0
3    253    0    0    0
3    212    0    0    0
3    201    0    0    0
3    179    0    0    0
3    186    0    0    0
3    198    0    0    0
3    244    0    0    0
3    193    0    0    0
3    249    0    0    0
3    209    0    0    0
3    272    0    0    0
3    208    0    0    0
3    204    0    0    0
3    178    0    0    0
3    277    0    0    0
3    239    0    0    0
3    242    0    0    0
3    200    0    0    0
3    174    0    0    0
3    189    0    0    0
3    250    0    0    0
3    194    0    0    0
3    185    0    0    0
3    211    0    0    0
3    210    0    0    0
3    275    0    0    0
3    169    0    0    0
3    252    0    0    0
