1    1694    0    1    0
1    188    0    1    0
1    191    0    1    0
1    265    0    1    0
1    1691    0    1    0
1    234    0    1    0
1    34    0    1    0
1    341    0    1    0
1    323    0    1    0
1    3717    0    1    0
1    109    0    1    0
1    24    0    1    0
1    280    0    1    0
1    126    0    1    0
1    88    0    1    0
1    468    0    1    0
1    264    0    1    0
1    348    0    1    0
1    118    0    1    0
1    3724    0    1    0
1    64    0    1    0
1    20    0    1    0
1    27    0    1    0
1    4115    0    1    0
1    131    0    1    0
1    164    0    1    0
1    273    0    1    0
1    122    0    1    0
1    411    0    1    0
1    3552    0    1    0
1    203    0    1    0
1    479    0    1    0
1    3548    0    1    0
1    226    0    1    0
1    556    0    1    0
1    3546    0    1    0
1    81    0    1    0
1    422    0    1    0
1    299    0    1    0
1    91    0    1    0
1    4090    0    1    0
1    52    0    1    0
1    26    0    1    0
1    315    0    1    0
1    112    0    1    0
1    167    0    1    0
1    386    0    1    0
1    332    0    1    0
1    1    0    1    0
1    136    0    1    0
1    23    0    1    0
1    4089    0    1    0
1    149    0    1    0
1    46    0    1    0
1    335    0    1    0
1    302    0    1    0
1    117    0    1    0
1    374    0    1    0
1    140    0    1    0
1    331    0    1    0
1    3550    0    1    0
1    158    0    1    0
1    257    0    1    0
1    137    0    1    0
1    549    0    1    0
1    87    0    1    0
1    113    0    1    0
1    173    0    1    0
1    176    0    1    0
1    70    0    1    0
1    435    0    1    0
1    490    0    1    0
1    103    0    1    0
1    86    0    1    0
1    245    0    1    0
1    141    0    1    0
1    80    0    1    0
1    94    0    1    0
1    31    0    1    0
1    248    0    1    0
1    218    0    1    0
1    1497    0    1    0
1    324    0    1    0
1    503    0    1    0
1    67    0    1    0
1    146    0    1    0
1    251    0    1    0
1    254    0    1    0
1    366    0    1    0
1    25    0    1    0
1    197    0    1    0
1    206    0    1    0
1    100    0    1    0
1    127    0    1    0
1    43    0    1    0
1    54    0    1    0
1    307    0    1    0
1    372    0    1    0
1    76    0    1    0
1    11    0    1    0
1    73    0    1    0
1    152    0    1    0
1    1689    0    1    0
1    97    0    1    0
1    2358    0    1    0
1    292    0    1    0
1    17    0    1    0
1    338    0    1    0
1    233    0    1    0
1    135    0    1    0
1    308    0    1    0
1    562    0    1    0
1    2174    0    1    0
1    145    0    1    0
1    400    0    1    0
1    182    0    1    0
1    225    0    1    0
1    79    0    1    0
1    241    0    1    0
1    61    0    1    0
1    373    0    1    0
1    4088    0    1    0
1    389    0    1    0
1    1690    0    1    0
1    53    0    1    0
1    4087    0    1    0
1    534    0    1    0
1    83    0    1    0
1    119    0    1    0
1    161    0    1    0
1    129    0    1    0
1    115    0    1    0
1    116    0    1    0
1    123    0    1    0
1    369    0    1    0
1    457    0    1    0
1    40    0    1    0
1    114    0    1    0
1    179    0    1    0
1    132    0    1    0
1    3173    0    1    0
1    293    0    1    0
1    281    0    1    0
1    288    0    1    0
1    4092    0    1    0
1    361    0    1    0
1    209    0    1    0
1    272    0    1    0
1    514    0    1    0
1    2824    0    1    0
1    289    0    1    0
1    316    0    1    0
1    559    0    1    0
1    82    0    1    0
1    170    0    1    0
1    4    0    1    0
1    120    0    1    0
1    106    0    1    0
1    14    0    1    0
1    130    0    1    0
1    446    0    1    0
1    242    0    1    0
1    200    0    1    0
1    351    0    1    0
1    37    0    1    0
1    358    0    1    0
1    552    0    1    0
1    4091    0    1    0
1    194    0    1    0
1    185    0    1    0
1    523    0    1    0
1    545    0    1    0
1    210    0    1    0
1    155    0    1    0
1    49    0    1    0
1    121    0    1    0
1    217    0    1    0
1    128    0    1    0
3    144    1    0    1    141
3    298    1    0    1    293
0    4114    7    1    2    135    4115
0    2825    5    1    1    2824
3    973    1    0    1    3173
0    3547    5    12    1    3546
0    3549    5    11    1    3548
0    3551    5    11    1    3550
0    3553    5    12    1    3552
3    594    5    0    1    545
3    599    5    0    1    348
3    600    5    0    1    366
3    601    7    0    2    552    562
3    602    5    0    1    549
3    603    5    0    1    545
3    604    5    0    1    545
3    611    5    0    1    338
3    612    5    0    1    358
0    633    6    1    2    373    1
3    810    7    0    2    141    145
0    814    5    1    1    3173
0    816    5    1    1    4114
0    844    7    1    2    2825    27
0    846    7    1    2    386    556
3    848    5    0    1    245
3    849    5    0    1    552
3    850    5    0    1    562
3    851    5    0    1    559
0    852    7    1    4    386    559    556    552
0    1502    5    3    1    1497
2    1528    1    1689
2    1552    1    1690
2    1609    1    1689
2    1633    1    1690
2    1697    1    137
2    1698    1    137
2    1701    1    141
0    2179    5    3    1    2174
2    2203    1    1691
2    2226    1    1694
2    2281    1    1691
2    2304    1    1694
2    2361    1    254
2    2370    1    251
2    2382    1    251
2    2393    1    248
2    2405    1    248
2    2418    1    4088
2    2442    1    4087
2    2476    1    4089
2    2500    1    4090
2    2533    1    210
2    2537    1    210
2    2541    1    218
2    2545    1    218
2    2549    1    226
2    2553    1    226
2    2557    1    234
2    2561    1    234
2    2627    1    257
2    2631    1    257
2    2635    1    265
2    2639    1    265
2    2643    1    273
2    2647    1    273
2    2651    1    281
2    2655    1    281
2    2721    1    335
2    2734    1    335
2    2816    1    206
0    2822    7    3    2    27    31
2    2826    1    1
2    2828    1    2358
2    2882    1    293
2    2886    1    302
2    2890    1    308
2    2894    1    308
2    2898    1    316
2    2902    1    316
2    2948    1    324
2    2952    1    324
2    2956    1    341
2    2960    1    341
2    2964    1    351
2    2968    1    351
2    3024    1    257
2    3028    1    257
2    3032    1    265
2    3036    1    265
2    3040    1    273
2    3044    1    273
2    3048    1    281
2    3052    1    281
2    3092    1    332
2    3105    1    332
2    3175    1    549
0    3176    7    4    2    31    27
0    3181    5    5    1    2358
2    3204    1    324
2    3208    1    324
2    3212    1    341
2    3216    1    341
2    3220    1    351
2    3224    1    351
2    3256    1    293
2    3260    1    302
2    3264    1    308
2    3268    1    308
2    3272    1    316
2    3276    1    316
2    3302    1    361
2    3314    1    361
2    3354    1    210
2    3358    1    210
2    3362    1    218
2    3366    1    218
2    3370    1    226
2    3374    1    226
2    3378    1    234
2    3382    1    234
0    3440    5    2    1    324
2    3554    1    242
2    3555    1    242
2    3556    1    254
2    3558    1    4088
2    3582    1    4087
2    3616    1    4092
2    3628    1    4091
2    3660    1    4089
2    3684    1    4090
0    3721    5    2    1    3717
0    3728    5    2    1    3724
2    3737    1    4091
2    3757    1    4092
2    3795    1    4091
2    3815    1    4092
2    3972    1    4091
2    3991    1    4092
2    4030    1    4091
2    4049    1    4092
2    4110    1    299
2    4119    1    446
2    4127    1    457
2    4135    1    468
2    4143    1    422
2    4151    1    435
2    4159    1    389
2    4167    1    400
2    4175    1    411
2    4183    1    374
2    4188    1    4
2    4276    1    446
2    4284    1    457
2    4292    1    468
2    4300    1    435
2    4308    1    389
2    4316    1    400
2    4324    1    411
2    4332    1    422
2    4340    1    374
2    4631    1    479
2    4639    1    490
2    4647    1    503
2    4655    1    514
2    4663    1    523
2    4671    1    534
2    4676    1    54
2    4764    1    479
2    4772    1    503
2    4780    1    514
2    4788    1    523
2    4796    1    534
2    4804    1    490
2    5082    1    361
2    5085    1    369
2    5090    1    341
2    5093    1    351
2    5098    1    308
2    5101    1    316
2    5108    1    293
2    5111    1    302
2    5332    1    281
2    5335    1    289
2    5340    1    265
2    5343    1    273
2    5348    1    234
2    5351    1    257
2    5356    1    218
2    5359    1    226
2    5369    1    210
3    634    5    0    1    633
3    815    7    0    2    136    814
3    845    5    0    1    844
3    847    5    0    1    846
3    926    1    0    1    1697
3    923    1    0    1    1701
3    921    1    0    1    2826
0    2979    7    1    2    3553    514
0    2999    3    1    2    3547    514
3    892    1    0    1    3175
3    887    1    0    1    4110
3    606    5    0    1    3175
0    1580    7    1    3    170    1528    1552
0    1586    7    1    3    173    1528    1552
0    1592    7    1    3    167    1528    1552
0    1598    7    1    3    164    1528    1552
0    1604    7    1    3    161    1528    1552
3    656    6    0    2    2822    140
0    1668    7    1    3    185    1609    1633
0    1674    7    1    3    158    1609    1633
0    1680    7    1    3    152    1609    1633
0    1686    7    1    3    146    1609    1633
0    2254    7    1    3    170    2203    2226
0    2260    7    1    3    173    2203    2226
0    2266    7    1    3    167    2203    2226
0    2272    7    1    3    164    2203    2226
0    2278    7    1    3    161    2203    2226
0    2339    7    1    3    185    2281    2304
0    2345    7    1    3    158    2281    2304
0    2351    7    1    3    152    2281    2304
0    2357    7    1    3    146    2281    2304
0    711    7    1    3    106    3660    3684
0    721    7    1    3    61    2418    2442
0    726    7    1    3    106    3558    3582
0    731    7    1    3    49    3558    3582
0    736    7    1    3    103    3558    3582
0    741    7    1    3    40    3558    3582
0    746    7    1    3    37    3558    3582
0    751    7    1    3    20    2418    2442
0    756    7    1    3    17    2418    2442
0    761    7    1    3    70    2418    2442
0    766    7    1    3    64    2418    2442
0    771    7    1    3    49    3660    3684
0    776    7    1    3    103    3660    3684
0    781    7    1    3    40    3660    3684
0    786    7    1    3    37    3660    3684
0    791    7    1    3    20    2476    2500
0    796    7    1    3    17    2476    2500
0    801    7    1    3    70    2476    2500
0    806    7    1    3    64    2476    2500
3    809    5    0    1    2822
0    3734    7    1    3    123    3728    3717
0    842    7    1    2    3795    3815
0    858    7    1    3    61    2476    2500
0    881    7    1    2    3737    3757
0    4123    5    1    1    4119
0    4131    5    1    1    4127
0    4139    5    1    1    4135
0    4147    5    1    1    4143
0    4155    5    1    1    4151
0    4163    5    1    1    4159
0    4171    5    1    1    4167
0    4179    5    1    1    4175
0    4187    5    1    1    4183
0    4194    5    1    1    4188
0    4282    5    1    1    4276
0    4290    5    1    1    4284
0    4298    5    1    1    4292
0    4306    5    1    1    4300
0    4314    5    1    1    4308
0    4322    5    1    1    4316
0    4330    5    1    1    4324
0    4338    5    1    1    4332
0    4346    5    1    1    4340
2    1526    1    1697
0    1540    5    10    1    1528
0    1564    5    10    1    1552
2    1606    1    1697
0    1621    5    10    1    1609
0    1645    5    10    1    1633
0    1661    7    1    3    179    1609    1633
2    1688    1    2826
0    4635    5    1    1    4631
0    4643    5    1    1    4639
0    4651    5    1    1    4647
0    4659    5    1    1    4655
0    4667    5    1    1    4663
0    4675    5    1    1    4671
0    4682    5    1    1    4676
0    4770    5    1    1    4764
0    4778    5    1    1    4772
0    4786    5    1    1    4780
0    4794    5    1    1    4788
0    4802    5    1    1    4796
0    4810    5    1    1    4804
2    2202    1    1698
0    2215    5    10    1    2203
0    2238    5    10    1    2226
2    2279    1    1698
0    2293    5    10    1    2281
0    2316    5    10    1    2304
0    2332    7    1    3    179    2281    2304
0    2430    5    10    1    2418
0    2454    5    10    1    2442
0    2488    5    10    1    2476
0    2512    5    10    1    2500
0    2536    5    1    1    2533
0    2540    5    1    1    2537
0    2544    5    1    1    2541
0    2548    5    1    1    2545
0    2552    5    1    1    2549
0    2556    5    1    1    2553
0    2560    5    1    1    2557
0    2564    5    1    1    2561
0    2566    7    1    3    3553    457    2537
0    2572    7    1    3    3553    468    2545
0    2578    7    1    3    3553    422    2553
0    2584    7    1    3    3553    435    2561
0    2590    7    1    2    3547    2533
0    2595    7    1    2    3547    2541
0    2600    7    1    2    3547    2549
0    2605    7    1    2    3547    2557
0    2630    5    1    1    2627
0    2634    5    1    1    2631
0    2638    5    1    1    2635
0    2642    5    1    1    2639
0    2646    5    1    1    2643
0    2650    5    1    1    2647
0    2654    5    1    1    2651
0    2658    5    1    1    2655
0    2660    7    1    3    3553    389    2631
0    2666    7    1    3    3553    400    2639
0    2672    7    1    3    3553    411    2647
0    2678    7    1    3    3553    374    2655
0    2684    7    1    2    3547    2627
0    2689    7    1    2    3547    2635
0    2694    7    1    2    3547    2643
0    2699    7    1    2    3547    2651
0    2728    5    5    1    2721
0    2741    5    5    1    2734
0    2748    7    1    2    292    2721
0    2750    7    1    2    288    2721
0    2752    7    1    2    280    2721
0    2754    7    1    2    272    2721
0    2756    7    1    2    264    2721
0    2758    7    1    2    241    2734
0    2760    7    1    2    233    2734
0    2762    7    1    2    225    2734
0    2764    7    1    2    217    2734
0    2766    7    1    2    209    2734
2    2827    1    1701
0    2838    5    8    1    2828
0    2847    5    9    1    2822
0    2885    5    1    1    2882
0    2889    5    1    1    2886
0    2893    5    1    1    2890
0    2897    5    1    1    2894
0    2901    5    1    1    2898
0    2905    5    1    1    2902
0    2906    7    1    2    2393    2886
0    2909    7    1    3    2393    479    2894
0    2913    7    1    3    2393    490    2902
0    2918    7    1    2    3554    2882
0    2922    7    1    2    3554    2890
0    2927    7    1    2    3554    2898
0    2951    5    1    1    2948
0    2955    5    1    1    2952
0    2959    5    1    1    2956
0    2963    5    1    1    2960
0    2967    5    1    1    2964
0    2971    5    1    1    2968
0    2973    7    1    3    3553    503    2952
0    2980    5    1    1    2979
0    2982    7    1    3    3553    523    2960
0    2988    7    1    3    3553    534    2968
0    2994    7    1    2    3547    2948
0    3001    7    1    2    3547    2956
0    3006    7    1    2    3547    2964
0    3027    5    1    1    3024
0    3031    5    1    1    3028
0    3035    5    1    1    3032
0    3039    5    1    1    3036
0    3043    5    1    1    3040
0    3047    5    1    1    3044
0    3051    5    1    1    3048
0    3055    5    1    1    3052
0    3056    7    1    3    2393    389    3028
0    3060    7    1    3    2393    400    3036
0    3064    7    1    3    2393    411    3044
0    3068    7    1    3    2393    374    3052
0    3073    7    1    2    3554    3024
0    3078    7    1    2    3554    3032
0    3083    7    1    2    3554    3040
0    3088    7    1    2    3554    3048
0    3099    5    5    1    3092
0    3112    5    5    1    3105
0    3119    7    1    2    372    3092
0    3121    7    1    2    366    3092
0    3123    7    1    2    358    3092
0    3125    7    1    2    348    3092
0    3126    7    1    2    338    3092
0    3128    7    1    2    331    3105
0    3130    7    1    2    323    3105
0    3132    7    1    2    315    3105
0    3134    7    1    2    307    3105
0    3136    7    1    2    299    3105
0    3187    5    4    1    3181
0    3193    7    1    2    83    3181
0    3196    7    1    2    86    3181
0    3199    7    1    2    88    3181
0    3202    7    1    2    88    3181
0    3207    5    1    1    3204
0    3211    5    1    1    3208
0    3215    5    1    1    3212
0    3219    5    1    1    3216
0    3223    5    1    1    3220
0    3227    5    1    1    3224
0    3228    7    1    3    2405    503    3208
0    3232    7    1    2    2405    514
0    3234    7    1    3    2405    523    3216
0    3238    7    1    3    2405    534    3224
0    3243    7    1    2    3555    3204
0    3247    3    1    2    3555    514
0    3249    7    1    2    3555    3212
0    3253    7    1    2    3555    3220
0    3259    5    1    1    3256
0    3263    5    1    1    3260
0    3267    5    1    1    3264
0    3271    5    1    1    3268
0    3275    5    1    1    3272
0    3279    5    1    1    3276
0    3280    7    1    2    2405    3260
0    3283    7    1    3    2405    479    3268
0    3287    7    1    3    2405    490    3276
0    3292    7    1    2    3555    3256
0    3295    7    1    2    3555    3264
0    3299    7    1    2    3555    3272
0    3305    5    1    1    3302
2    3306    1    2816
2    3310    1    2816
0    3317    5    1    1    3314
2    3318    1    2816
2    3322    1    2816
0    3326    7    1    2    2405    3302
0    3333    7    1    2    2405    3314
0    3357    5    1    1    3354
0    3361    5    1    1    3358
0    3365    5    1    1    3362
0    3369    5    1    1    3366
0    3373    5    1    1    3370
0    3377    5    1    1    3374
0    3381    5    1    1    3378
0    3385    5    1    1    3382
0    3386    7    1    3    2393    457    3358
0    3390    7    1    3    2393    468    3366
0    3394    7    1    3    2393    422    3374
0    3398    7    1    3    2393    435    3382
0    3403    7    1    2    3554    3354
0    3408    7    1    2    3554    3362
0    3413    7    1    2    3554    3370
0    3418    7    1    2    3554    3378
0    5088    5    1    1    5082
0    5089    5    1    1    5085
0    5096    5    1    1    5090
0    5097    5    1    1    5093
2    3489    1    3440
2    3493    1    3440
0    3570    5    10    1    3558
0    3594    5    10    1    3582
0    3622    5    4    1    3616
0    3632    5    2    1    3628
0    3637    7    1    2    97    3616
0    3640    7    1    2    94    3616
0    3643    7    1    2    97    3616
0    3646    7    1    2    94    3616
0    3672    5    10    1    3660
0    3696    5    10    1    3684
0    3745    5    10    1    3737
0    3765    5    10    1    3757
0    3803    5    10    1    3795
0    3823    5    10    1    3815
0    5338    5    1    1    5332
0    5339    5    1    1    5335
0    5346    5    1    1    5340
0    5347    5    1    1    5343
0    5354    5    1    1    5348
0    5355    5    1    1    5351
0    3979    5    10    1    3972
0    3998    5    10    1    3991
0    4037    5    10    1    4030
0    4056    5    10    1    4049
2    4094    1    4110
0    5104    5    1    1    5098
0    5105    5    1    1    5101
0    5114    5    1    1    5108
0    5115    5    1    1    5111
0    5362    5    1    1    5356
0    5363    5    1    1    5359
2    5366    1    2816
0    5373    5    1    1    5369
3    993    1    0    1    1688
3    978    1    0    1    1688
3    949    1    0    1    1688
3    939    1    0    1    1688
0    2568    7    1    3    457    3551    2540
0    2574    7    1    3    468    3551    2548
0    2580    7    1    3    422    3551    2556
0    2586    7    1    3    435    3551    2564
0    2592    7    1    2    3549    2536
0    2597    7    1    2    3549    2544
0    2602    7    1    2    3549    2552
0    2607    7    1    2    3549    2560
0    2662    7    1    3    389    3551    2634
0    2668    7    1    3    400    3551    2642
0    2674    7    1    3    411    3551    2650
0    2680    7    1    3    374    3551    2658
0    2686    7    1    2    3549    2630
0    2691    7    1    2    3549    2638
0    2696    7    1    2    3549    2646
0    2701    7    1    2    3549    2654
0    2907    7    1    2    2370    2889
0    2910    7    1    3    479    2370    2897
0    2914    7    1    3    490    2370    2905
0    2920    7    1    2    3556    2885
0    2924    7    1    2    3556    2893
0    2929    7    1    2    3556    2901
0    2975    7    1    3    503    3551    2955
0    2984    7    1    3    523    3551    2963
0    2990    7    1    3    534    3551    2971
0    2996    7    1    2    3549    2951
0    3003    7    1    2    3549    2959
0    3008    7    1    2    3549    2967
0    3015    7    2    2    2980    2999
0    3057    7    1    3    389    2370    3031
0    3061    7    1    3    400    2370    3039
0    3065    7    1    3    411    2370    3047
0    3069    7    1    3    374    2370    3055
0    3075    7    1    2    3556    3027
0    3080    7    1    2    3556    3035
0    3085    7    1    2    3556    3043
0    3090    7    1    2    3556    3051
0    3229    7    1    3    503    2382    3211
0    3233    5    1    1    3232
0    3235    7    1    3    523    2382    3219
0    3239    7    1    3    534    2382    3227
0    3244    7    1    2    2361    3207
0    3250    7    1    2    2361    3215
0    3254    7    1    2    2361    3223
0    3281    7    1    2    2382    3263
0    3284    7    1    3    479    2382    3271
0    3288    7    1    3    490    2382    3279
0    3293    7    1    2    2361    3259
0    3296    7    1    2    2361    3267
0    3300    7    1    2    2361    3275
0    3327    7    1    2    2382    3305
0    3334    7    1    2    2382    3317
0    3387    7    1    3    457    2370    3361
0    3391    7    1    3    468    2370    3369
0    3395    7    1    3    422    2370    3377
0    3399    7    1    3    435    2370    3385
0    3405    7    1    2    3556    3357
0    3410    7    1    2    3556    3365
0    3415    7    1    2    3556    3373
0    3420    7    1    2    3556    3381
0    3422    6    1    2    5085    5088
0    3423    6    1    2    5082    5089
0    3431    6    1    2    5093    5096
0    3432    6    1    2    5090    5097
0    3895    6    1    2    5335    5338
0    3896    6    1    2    5332    5339
0    3904    6    1    2    5343    5346
0    3905    6    1    2    5340    5347
0    3913    6    1    2    5351    5354
0    3914    6    1    2    5348    5355
3    889    1    0    1    4094
0    5106    6    1    2    5101    5104
0    5107    6    1    2    5098    5105
0    5116    6    1    2    5111    5114
0    5117    6    1    2    5108    5115
0    5364    6    1    2    5359    5362
0    5365    6    1    2    5356    5363
3    593    5    0    1    4094
0    2880    7    1    2    2838    2847
0    2881    7    1    2    2828    2847
0    1579    7    1    3    200    1540    1552
0    1585    7    1    3    203    1540    1552
0    1591    7    1    3    197    1540    1552
0    1597    7    1    3    194    1540    1552
0    1603    7    1    3    191    1540    1552
0    1667    7    1    3    182    1621    1633
0    1673    7    1    3    188    1621    1633
0    1679    7    1    3    155    1621    1633
0    1685    7    1    3    149    1621    1633
0    2876    7    1    2    2838    2847
0    2877    7    1    2    2828    2847
0    2253    7    1    3    200    2215    2226
0    2259    7    1    3    203    2215    2226
0    2265    7    1    3    197    2215    2226
0    2271    7    1    3    194    2215    2226
0    2277    7    1    3    191    2215    2226
0    2338    7    1    3    182    2293    2304
0    2344    7    1    3    188    2293    2304
0    2350    7    1    3    155    2293    2304
0    2356    7    1    3    149    2293    2304
0    2868    7    1    2    2838    2847
0    2869    7    1    2    2828    2847
0    710    7    1    3    109    3672    3684
0    2872    7    1    2    2838    2847
0    2873    7    1    2    2828    2847
0    720    7    1    3    11    2430    2442
0    725    7    1    3    109    3570    3582
0    730    7    1    3    46    3570    3582
0    735    7    1    3    100    3570    3582
0    740    7    1    3    91    3570    3582
0    745    7    1    3    43    3570    3582
0    750    7    1    3    76    2430    2442
0    755    7    1    3    73    2430    2442
0    760    7    1    3    67    2430    2442
0    765    7    1    3    14    2430    2442
0    770    7    1    3    46    3672    3684
0    775    7    1    3    100    3672    3684
0    780    7    1    3    91    3672    3684
0    785    7    1    3    43    3672    3684
0    790    7    1    3    76    2488    2500
0    795    7    1    3    73    2488    2500
0    800    7    1    3    67    2488    2500
0    805    7    1    3    14    2488    2500
0    841    7    1    3    120    3803    3815
0    857    7    1    3    11    2488    2500
0    880    7    1    3    118    3745    3757
0    1660    7    1    3    176    1621    1633
0    2331    7    1    3    176    2293    2304
0    2569    3    1    2    2566    2568
0    2575    3    1    2    2572    2574
0    2581    3    1    2    2578    2580
0    2587    3    1    2    2584    2586
0    2593    3    1    3    2590    2592    457
0    2598    3    1    3    2595    2597    468
0    2603    3    1    3    2600    2602    422
0    2608    3    1    3    2605    2607    435
0    2663    3    1    2    2660    2662
0    2669    3    1    2    2666    2668
0    2675    3    1    2    2672    2674
0    2681    3    1    2    2678    2680
0    2687    3    1    3    2684    2686    389
0    2692    3    1    3    2689    2691    400
0    2697    3    1    3    2694    2696    411
0    2702    3    1    3    2699    2701    374
0    2747    7    1    2    289    2728
0    2749    7    1    2    281    2728
0    2751    7    1    2    273    2728
0    2753    7    1    2    265    2728
0    2755    7    1    2    257    2728
0    2757    7    1    2    234    2741
0    2759    7    1    2    226    2741
0    2761    7    1    2    218    2741
0    2763    7    1    2    210    2741
0    2765    7    1    2    206    2741
0    2857    5    8    1    2847
0    2908    3    1    2    2906    2907
0    2911    3    1    2    2909    2910
0    2915    3    1    2    2913    2914
0    2925    3    1    3    2922    2924    479
0    2930    3    1    3    2927    2929    490
0    2933    3    2    2    2918    2920
0    2976    3    1    2    2973    2975
0    2985    3    1    2    2982    2984
0    2991    3    1    2    2988    2990
0    2997    3    1    3    2994    2996    503
0    3004    3    1    3    3001    3003    523
0    3009    3    1    3    3006    3008    534
0    3058    3    1    2    3056    3057
0    3062    3    1    2    3060    3061
0    3066    3    1    2    3064    3065
0    3070    3    1    2    3068    3069
0    3076    3    1    3    3073    3075    389
0    3081    3    1    3    3078    3080    400
0    3086    3    1    3    3083    3085    411
0    3091    3    1    3    3088    3090    374
0    3118    7    1    2    369    3099
0    3120    7    1    2    361    3099
0    3122    7    1    2    351    3099
0    3124    7    1    2    341    3099
0    3127    7    1    2    324    3112
0    3129    7    1    2    316    3112
0    3131    7    1    2    308    3112
0    3133    7    1    2    302    3112
0    3135    7    1    2    293    3112
0    3147    3    5    2    3099    3126
0    3192    7    1    2    83    3187
0    3195    7    1    2    87    3187
0    3198    7    1    2    34    3187
0    3201    7    1    2    34    3187
0    3230    3    1    2    3228    3229
0    3236    3    1    2    3234    3235
0    3240    3    1    2    3238    3239
0    3245    3    1    3    3243    3244    503
0    3251    3    1    3    3249    3250    523
0    3255    3    1    3    3253    3254    534
0    3282    3    1    2    3280    3281
0    3285    3    1    2    3283    3284
0    3289    3    1    2    3287    3288
0    3297    3    1    3    3295    3296    479
0    3301    3    1    3    3299    3300    490
0    3309    5    1    1    3306
0    3313    5    1    1    3310
0    3321    5    1    1    3318
0    3325    5    1    1    3322
0    3328    3    1    2    3326    3327
0    3329    7    1    3    2405    446    3310
0    3335    3    1    2    3333    3334
0    3336    7    1    3    2405    446    3322
0    3341    7    1    2    3555    3306
0    3345    7    1    2    3555    3318
0    3388    3    1    2    3386    3387
0    3392    3    1    2    3390    3391
0    3396    3    1    2    3394    3395
0    3400    3    1    2    3398    3399
0    3406    3    1    3    3403    3405    457
0    3411    3    1    3    3408    3410    468
0    3416    3    1    3    3413    3415    422
0    3421    3    1    3    3418    3420    435
0    3424    6    3    2    3422    3423
0    3433    6    3    2    3431    3432
0    3492    5    1    1    3489
0    3496    5    1    1    3493
0    3780    7    1    3    117    3745    3757
0    3783    7    1    3    126    3745    3757
0    3786    7    1    3    127    3745    3757
0    3789    7    1    3    128    3745    3757
0    3838    7    1    3    131    3803    3815
0    3841    7    1    3    129    3803    3815
0    3844    7    1    3    119    3803    3815
0    3847    7    1    3    130    3803    3815
0    3897    6    3    2    3895    3896
0    3906    6    3    2    3904    3905
0    3915    6    2    2    3913    3914
0    4011    7    1    3    122    3979    3991
0    4014    7    1    3    113    3979    3991
0    4017    7    1    3    53    3979    3991
0    4020    7    1    3    114    3979    3991
0    4023    7    1    3    115    3979    3991
0    4069    7    1    3    52    4037    4049
0    4072    7    1    3    112    4037    4049
0    4075    7    1    3    116    4037    4049
0    4078    7    1    3    121    4037    4049
0    4081    7    1    3    123    4037    4049
0    5206    6    2    2    5116    5117
0    5209    6    2    2    5106    5107
0    5307    7    2    2    3233    3247
0    5322    3    2    2    3292    3293
0    5372    5    1    1    5366
0    5375    6    1    2    5366    5373
0    5399    6    2    2    5364    5365
0    2813    5    1    1    3015
0    3197    3    1    2    3195    3196
0    3200    3    1    2    3198    3199
0    3203    3    1    2    3201    3202
0    3194    3    1    2    3192    3193
0    2570    5    1    1    2569
0    2576    5    1    1    2575
0    2582    5    1    1    2581
0    2588    5    1    1    2587
0    2664    5    1    1    2663
0    2670    5    1    1    2669
0    2676    5    1    1    2675
0    2682    5    1    1    2681
0    2767    3    6    2    2749    2750
0    2772    3    5    2    2751    2752
0    2776    3    5    2    2753    2754
0    2780    3    5    2    2755    2756
0    2784    3    5    2    2757    2758
0    2788    3    7    2    2759    2760
0    2794    3    5    2    2761    2762
0    2798    3    5    2    2763    2764
0    2802    3    5    2    2765    2766
0    2912    5    1    1    2911
0    2916    5    1    1    2915
0    2936    5    2    1    2908
0    2977    5    1    1    2976
0    2986    5    1    1    2985
0    2992    5    1    1    2991
0    3059    5    1    1    3058
0    3063    5    1    1    3062
0    3067    5    1    1    3066
0    3071    5    1    1    3070
0    3137    3    5    2    3120    3121
0    3139    3    5    2    3122    3123
0    3143    3    5    2    3124    3125
0    3151    3    5    2    3127    3128
0    3155    3    7    2    3129    3130
0    3161    3    5    2    3131    3132
0    3165    3    5    2    3133    3134
0    3167    3    6    2    3135    3136
0    3231    5    1    1    3230
0    3237    5    1    1    3236
0    3241    5    1    1    3240
0    3286    5    1    1    3285
0    3290    5    1    1    3289
0    3330    7    1    3    446    2382    3313
0    3337    7    1    3    446    2382    3325
0    3342    7    1    2    2361    3309
0    3346    7    1    2    2361    3321
0    3348    5    2    1    3328
0    3352    5    1    1    3335
0    3389    5    1    1    3388
0    3393    5    1    1    3392
0    3397    5    1    1    3396
0    3401    5    1    1    3400
0    3845    7    1    3    3015    3803    3823
0    5126    3    2    2    3118    3119
0    5178    3    2    2    2747    2748
0    5325    5    2    1    3282
0    5374    6    1    2    5369    5372
0    2810    5    1    1    2933
0    635    7    1    2    3197    3176
0    2878    7    1    3    24    2838    2857
0    2879    7    1    3    25    2828    2857
0    2874    7    1    3    26    2838    2857
0    2875    7    1    3    81    2828    2857
0    703    7    1    2    3200    3176
0    2866    7    1    3    79    2838    2857
0    2867    7    1    3    23    2828    2857
0    2870    7    1    3    82    2838    2857
0    2871    7    1    3    80    2828    2857
0    716    7    1    2    3203    3176
0    819    7    1    2    3194    3176
0    1789    7    2    2    3147    514
0    2036    7    3    2    514    3147
0    2611    7    2    2    2570    2593
0    2615    7    2    2    2576    2598
0    2619    7    2    2    2582    2603
0    2623    7    2    2    2588    2608
0    2705    7    2    2    2664    2687
0    2709    7    2    2    2670    2692
0    2713    7    2    2    2676    2697
0    2717    7    2    2    2682    2702
0    2939    7    2    2    2912    2925
0    2942    7    2    2    2916    2930
2    2945    1    2933
0    3012    7    2    2    2977    2997
0    3018    7    2    2    2986    3004
0    3021    7    2    2    2992    3009
0    3331    3    1    2    3329    3330
0    3338    3    1    2    3336    3337
0    3343    3    1    3    3341    3342    446
0    3347    3    1    3    3345    3346    446
0    3428    5    2    1    3424
0    3437    5    2    1    3433
0    3514    7    1    3    3433    3424    3489
0    3836    7    1    3    3352    3803    3823
0    3852    7    1    2    3071    3091
0    5311    5    1    1    5307
0    3901    5    2    1    3897
0    3910    5    2    1    3906
2    3934    1    3915
2    3938    1    3915
2    4652    1    3147
2    4783    1    3147
2    5137    1    3147
0    5212    5    1    1    5206
0    5213    5    1    1    5209
0    5260    7    2    2    3063    3081
0    5263    7    2    2    3067    3086
0    5268    7    2    2    3401    3421
0    5271    7    2    2    3059    3076
0    5276    7    2    2    3393    3411
0    5279    7    2    2    3397    3416
0    5289    7    2    2    3389    3406
0    5296    7    2    2    3237    3251
0    5299    7    2    2    3241    3255
0    5304    7    2    2    3231    3245
0    5312    7    2    2    3286    3297
0    5315    7    2    2    3290    3301
0    5328    5    1    1    5322
0    5396    6    2    2    5374    5375
0    5403    5    1    1    5399
0    1286    7    1    2    446    2802
0    2809    5    1    1    2936
0    597    5    1    1    3348
0    1031    7    1    2    2802    446
3    636    5    0    1    635
0    637    3    1    4    2878    2879    2880    2881
0    671    3    1    4    2874    2875    2876    2877
3    704    5    0    1    703
0    705    3    1    4    2866    2867    2868    2869
0    713    3    1    4    2870    2871    2872    2873
3    717    5    0    1    716
3    820    5    0    1    819
0    1046    7    3    2    2798    457
0    1064    7    5    2    2794    468
0    1071    7    6    2    422    2788
0    1097    7    1    2    2784    435
0    1111    7    2    2    2780    389
0    1128    7    3    2    2776    400
0    1145    7    4    2    2772    411
0    1160    7    5    2    2767    374
0    1301    7    3    2    457    2798
0    1318    7    4    2    468    2794
0    1324    7    5    2    422    2788
0    1341    7    1    2    435    2784
0    1359    7    3    2    389    2780
0    1382    7    5    2    400    2776
0    1404    7    6    2    411    2772
0    1412    7    7    2    374    2767
0    1704    5    6    1    3167
0    1712    5    10    1    3165
2    1724    1    3165
0    1742    7    5    2    3161    479
0    1749    7    6    2    490    3155
0    1775    7    1    2    3151    503
0    1806    7    3    2    3143    523
0    1823    7    4    2    3139    534
0    1829    5    6    1    3137
2    1837    1    3137
0    1958    5    6    1    3167
0    1966    5    10    1    3165
2    1978    1    3165
0    1995    7    4    2    479    3161
0    2001    7    5    2    490    3155
0    2018    7    1    2    503    3151
0    2059    7    5    2    523    3143
0    2081    7    6    2    534    3139
2    2089    1    3137
0    2106    5    6    1    3137
2    3170    1    3167
0    3332    5    1    1    3331
0    3339    5    1    1    3338
0    5132    5    1    1    5126
0    5184    5    1    1    5178
0    3853    5    3    1    3852
0    3874    5    3    1    3348
0    4076    7    1    3    2936    4037    4056
2    4116    1    2802
2    4124    1    2798
2    4132    1    2794
2    4140    1    2788
2    4148    1    2784
2    4156    1    2780
2    4164    1    2776
2    4172    1    2772
2    4180    1    2767
0    4228    4    2    2    422    2788
2    4279    1    2802
2    4287    1    2798
2    4295    1    2794
2    4303    1    2784
2    4311    1    2780
2    4319    1    2776
2    4327    1    2772
2    4335    1    2788
2    4343    1    2767
0    4348    4    2    2    422    2788
0    4464    4    2    2    374    2767
2    4628    1    3161
2    4636    1    3155
2    4644    1    3151
2    4660    1    3143
2    4668    1    3139
0    4716    4    2    2    490    3155
2    4767    1    3161
2    4775    1    3151
2    4791    1    3143
2    4799    1    3139
2    4807    1    3155
0    4812    4    2    2    490    3155
2    5118    1    3139
2    5121    1    3143
2    5129    1    3137
2    5134    1    3151
2    5142    1    3161
2    5145    1    3155
2    5152    1    3167
2    5155    1    3165
2    5162    1    2788
2    5165    1    2784
2    5170    1    2798
2    5173    1    2794
2    5181    1    2802
2    5186    1    2772
2    5189    1    2767
2    5196    1    2780
2    5199    1    2776
0    5214    6    1    2    5209    5212
0    5215    6    1    2    5206    5213
0    5329    5    1    1    5325
0    5330    6    1    2    5325    5328
0    2807    5    1    1    2942
0    2808    5    1    1    2939
0    2811    5    1    1    3021
0    2812    5    1    1    3018
0    2814    5    1    1    3012
0    2626    5    1    1    2623
0    2622    5    1    1    2619
0    2618    5    1    1    2615
0    2614    5    1    1    2611
0    2720    5    1    1    2717
0    2716    5    1    1    2713
0    2712    5    1    1    2709
0    2708    5    1    1    2705
3    639    7    0    2    637    2827
3    673    7    0    2    671    2827
3    707    7    0    2    705    2827
3    715    7    0    2    713    2827
0    3731    7    1    3    2945    3728    3721
0    4658    5    1    1    4652
0    1777    6    1    2    4652    4659
0    2019    6    1    2    4783    4786
0    4787    5    1    1    4783
0    3350    7    2    2    3332    3343
0    3353    7    1    2    3339    3347
0    5141    5    1    1    5137
0    3513    7    1    3    3428    3433    3492
0    3516    7    1    3    3424    3437    3496
0    3517    7    1    3    3437    3428    3493
0    3778    7    1    3    2717    3745    3765
0    3781    7    1    3    2713    3745    3765
0    3784    7    1    3    2709    3745    3765
0    3787    7    1    3    2705    3745    3765
0    3839    7    1    3    3021    3803    3823
0    3842    7    1    3    3018    3803    3823
0    5266    5    1    1    5260
0    5267    5    1    1    5263
0    5274    5    1    1    5268
0    5275    5    1    1    5271
0    5302    5    1    1    5296
0    5303    5    1    1    5299
0    5310    5    1    1    5304
0    3891    6    1    2    5304    5311
0    3937    5    1    1    3934
0    3941    5    1    1    3938
0    3955    7    1    3    3906    3897    3934
0    3958    7    1    3    3910    3901    3938
0    4009    7    1    3    2623    3979    3998
0    4012    7    1    3    2619    3979    3998
0    4015    7    1    3    2615    3979    3998
0    4018    7    1    3    2611    3979    3998
0    4067    7    1    3    3012    4037    4056
0    4070    7    1    3    2942    4037    4056
0    4073    7    1    3    2939    4037    4056
0    4079    7    1    3    2945    4037    4056
0    5239    6    2    2    5214    5215
0    5282    5    1    1    5276
0    5283    5    1    1    5279
0    5293    5    1    1    5289
0    5318    5    1    1    5312
0    5319    5    1    1    5315
0    5331    6    1    2    5322    5329
0    5402    5    1    1    5396
0    5405    6    1    2    5396    5403
0    595    7    1    4    2807    2808    2809    2810
0    596    7    1    4    2811    2812    2813    2814
0    607    7    1    4    2626    2622    2618    2614
0    608    7    1    4    2720    2716    2712    2708
0    1845    7    1    2    1704    1724
0    1846    7    1    3    1712    1704    1742
0    2115    7    1    2    1958    1978
0    2116    7    1    3    1966    1958    1995
0    4122    5    1    1    4116
0    1022    6    1    2    4116    4123
0    4130    5    1    1    4124
0    1033    6    1    2    4124    4131
0    4138    5    1    1    4132
0    1051    6    1    2    4132    4139
0    4146    5    1    1    4140
0    1079    6    1    2    4140    4147
0    4154    5    1    1    4148
0    1088    6    1    2    4148    4155
0    4162    5    1    1    4156
0    1099    6    1    2    4156    4163
0    4170    5    1    1    4164
0    1115    6    1    2    4164    4171
0    4178    5    1    1    4172
0    1133    6    1    2    4172    4179
0    4186    5    1    1    4180
0    1151    6    1    2    4180    4187
0    4234    5    1    1    4228
0    1276    6    1    2    4279    4282
0    4283    5    1    1    4279
0    1287    6    1    2    4287    4290
0    4291    5    1    1    4287
0    1305    6    1    2    4295    4298
0    4299    5    1    1    4295
0    1330    6    1    2    4303    4306
0    4307    5    1    1    4303
0    1342    6    1    2    4311    4314
0    4315    5    1    1    4311
0    1363    6    1    2    4319    4322
0    4323    5    1    1    4319
0    1388    6    1    2    4327    4330
0    4331    5    1    1    4327
0    1420    6    1    2    4335    4338
0    4339    5    1    1    4335
0    1428    6    1    2    4343    4346
0    4347    5    1    1    4343
0    4634    5    1    1    4628
0    1729    6    1    2    4628    4635
0    4642    5    1    1    4636
0    1757    6    1    2    4636    4643
0    4650    5    1    1    4644
0    1766    6    1    2    4644    4651
0    1776    6    1    2    4655    4658
0    4666    5    1    1    4660
0    1793    6    1    2    4660    4667
0    4674    5    1    1    4668
0    1811    6    1    2    4668    4675
0    1849    7    1    2    1712    1742
0    1852    7    1    2    1712    1742
0    1875    7    1    2    54    1829
0    4722    5    1    1    4716
0    1982    6    1    2    4767    4770
0    4771    5    1    1    4767
0    2007    6    1    2    4775    4778
0    4779    5    1    1    4775
0    2020    6    1    2    4780    4787
0    2040    6    1    2    4791    4794
0    4795    5    1    1    4791
0    2065    6    1    2    4799    4802
0    4803    5    1    1    4799
0    2097    6    1    2    4807    4810
0    4811    5    1    1    4807
0    2119    7    1    2    1966    1995
0    2122    7    1    2    1966    1995
0    5124    5    1    1    5118
0    5125    5    1    1    5121
0    3452    6    1    2    5129    5132
0    5133    5    1    1    5129
0    5140    5    1    1    5134
0    3462    6    1    2    5134    5141
0    5168    5    1    1    5162
0    5169    5    1    1    5165
0    5176    5    1    1    5170
0    5177    5    1    1    5173
0    3484    6    1    2    5181    5184
0    5185    5    1    1    5181
0    3515    4    1    2    3513    3514
0    3518    4    1    2    3516    3517
0    3857    5    2    1    3853
0    3860    6    1    2    5263    5266
0    3861    6    1    2    5260    5267
0    3869    6    1    2    5271    5274
0    3870    6    1    2    5268    5275
0    3878    5    2    1    3874
0    3881    6    1    2    5299    5302
0    3882    6    1    2    5296    5303
0    3890    6    1    2    5307    5310
0    3954    7    1    3    3901    3906    3937
0    3957    7    1    3    3897    3910    3941
0    4021    7    1    3    3353    3979    3998
0    4099    5    2    1    3170
2    4236    1    1071
0    4354    5    1    1    4348
2    4406    1    1324
0    4470    5    1    1    4464
2    4552    1    1412
2    4679    1    1829
2    4687    1    1704
2    4695    1    1704
2    4703    1    1712
2    4711    1    1712
2    4724    1    1749
0    4818    5    1    1    4812
2    4855    1    1958
2    4865    1    1966
2    4870    1    2001
2    4913    1    1958
2    4923    1    1966
2    4951    1    2106
2    5006    1    2089
2    5039    1    2106
0    5148    5    1    1    5142
0    5149    5    1    1    5145
0    5158    5    1    1    5152
0    5159    5    1    1    5155
0    5192    5    1    1    5186
0    5193    5    1    1    5189
0    5202    5    1    1    5196
0    5203    5    1    1    5199
0    5284    6    1    2    5279    5282
0    5285    6    1    2    5276    5283
0    5320    6    1    2    5315    5318
0    5321    6    1    2    5312    5319
0    5386    6    2    2    5330    5331
0    5404    6    1    2    5399    5402
3    598    7    0    3    595    596    597
0    609    5    1    1    3350
0    1021    6    1    2    4119    4122
0    1032    6    1    2    4127    4130
0    1050    6    1    2    4135    4138
0    1078    6    1    2    4143    4146
0    1087    6    1    2    4151    4154
0    1098    6    1    2    4159    4162
0    1114    6    1    2    4167    4170
0    1132    6    1    2    4175    4178
0    1150    6    1    2    4183    4186
0    1277    6    1    2    4276    4283
0    1288    6    1    2    4284    4291
0    1306    6    1    2    4292    4299
0    1331    6    1    2    4300    4307
0    1343    6    1    2    4308    4315
0    1364    6    1    2    4316    4323
0    1389    6    1    2    4324    4331
0    1421    6    1    2    4332    4339
0    1429    6    1    2    4340    4347
0    1728    6    1    2    4631    4634
0    1756    6    1    2    4639    4642
0    1765    6    1    2    4647    4650
0    1778    6    9    2    1776    1777
0    1792    6    1    2    4663    4666
0    1810    6    1    2    4671    4674
0    1983    6    1    2    4764    4771
0    2008    6    1    2    4772    4779
0    2021    6    13    2    2019    2020
0    2041    6    1    2    4788    4795
0    2066    6    1    2    4796    4803
0    2098    6    1    2    4804    4811
0    3443    6    1    2    5121    5124
0    3444    6    1    2    5118    5125
0    3453    6    1    2    5126    5133
0    3461    6    1    2    5137    5140
0    3466    6    1    2    5165    5168
0    3467    6    1    2    5162    5169
0    3475    6    1    2    5173    5176
0    3476    6    1    2    5170    5177
0    3485    6    1    2    5178    5185
0    5243    5    1    1    5239
0    3862    6    3    2    3860    3861
0    3871    6    2    2    3869    3870
0    3883    6    3    2    3881    3882
0    3892    6    2    2    3890    3891
0    3956    4    1    2    3954    3955
0    3959    4    1    2    3957    3958
0    4756    3    2    2    1837    1875
0    5150    6    1    2    5145    5148
0    5151    6    1    2    5142    5149
0    5160    6    1    2    5155    5158
0    5161    6    1    2    5152    5159
0    5194    6    1    2    5189    5192
0    5195    6    1    2    5186    5193
0    5204    6    1    2    5199    5202
0    5205    6    1    2    5196    5203
0    5236    6    2    2    3518    3515
2    5286    1    3350
0    5379    6    2    2    5284    5285
0    5389    6    2    2    5320    5321
0    5425    6    2    2    5404    5405
3    610    7    0    3    607    608    609
0    1023    6    6    2    1021    1022
0    1034    6    10    2    1032    1033
0    1052    6    10    2    1050    1051
0    1080    6    5    2    1078    1079
0    1089    6    6    2    1087    1088
0    1100    6    9    2    1098    1099
0    1116    6    10    2    1114    1115
0    1134    6    9    2    1132    1133
0    1152    6    6    2    1150    1151
0    4242    5    1    1    4236
0    1278    6    6    2    1276    1277
0    1289    6    10    2    1287    1288
0    1307    6    9    2    1305    1306
0    1332    6    7    2    1330    1331
0    1344    6    13    2    1342    1343
0    1365    6    15    2    1363    1364
0    1390    6    12    2    1388    1389
0    1422    6    5    2    1420    1421
0    1430    6    6    2    1428    1429
0    1730    6    10    2    1728    1729
0    1758    6    5    2    1756    1757
0    1767    6    6    2    1765    1766
0    1794    6    10    2    1792    1793
0    1812    6    9    2    1810    1811
0    1876    6    1    2    4679    4682
0    4683    5    1    1    4679
0    4691    5    1    1    4687
0    4699    5    1    1    4695
0    4707    5    1    1    4703
0    4715    5    1    1    4711
0    4730    5    1    1    4724
0    1984    6    9    2    1982    1983
0    2009    6    7    2    2007    2008
0    2042    6    15    2    2040    2041
0    2067    6    12    2    2065    2066
0    2099    6    5    2    2097    2098
0    4869    5    1    1    4865
0    4927    5    1    1    4923
0    3445    6    3    2    3443    3444
0    3454    6    3    2    3452    3453
0    3463    6    2    2    3461    3462
0    3468    6    3    2    3466    3467
0    3477    6    3    2    3475    3476
0    3486    6    2    2    3484    3485
0    4103    7    1    2    4099    3170
0    4412    5    1    1    4406
0    4558    5    1    1    4552
0    4859    5    1    1    4855
0    4876    5    1    1    4870
0    4917    5    1    1    4913
0    4955    5    1    1    4951
0    5012    5    1    1    5006
0    5043    5    1    1    5039
0    5216    6    2    2    5160    5161
0    5219    6    2    2    5150    5151
0    5226    6    2    2    5204    5205
0    5229    6    2    2    5194    5195
0    5392    5    1    1    5386
0    5422    6    2    2    3959    3956
0    1866    7    1    2    1778    1806
0    1877    6    1    2    4676    4683
0    4762    5    1    1    4756
0    2142    7    1    2    2021    2059
0    2146    7    1    2    2021    2059
0    5242    5    1    1    5236
0    3532    6    1    2    5236    5243
0    3866    5    2    1    3862
0    3887    5    2    1    3883
2    3918    1    3871
2    3922    1    3871
2    3926    1    3892
2    3930    1    3892
0    5429    5    1    1    5425
0    4104    3    2    2    4099    4103
2    4743    1    1778
2    4991    1    2021
2    5001    1    2021
0    5292    5    1    1    5286
0    5295    6    1    2    5286    5293
0    5383    5    1    1    5379
0    5393    5    1    1    5389
0    5394    6    1    2    5389    5392
0    1439    7    1    2    1278    1301
0    1440    7    1    3    1289    1278    1318
0    1441    7    1    4    1307    1278    1324    1289
0    1847    7    1    4    1730    1704    1749    1712
0    1168    7    1    2    1023    1046
0    1169    7    1    3    1034    1023    1064
0    1170    7    1    4    1052    1023    1071    1034
0    2117    7    1    4    1984    1958    2001    1966
0    1086    5    1    1    1080
0    1166    7    2    4    1034    1080    1052    1023
0    1171    7    1    2    1034    1064
0    1172    7    1    3    1052    1071    1034
0    1173    7    1    3    1080    1052    1034
0    1174    7    1    2    1034    1064
0    1175    7    1    3    1071    1052    1034
0    1176    7    1    2    1052    1071
0    1177    7    1    2    1080    1052
0    1178    7    1    2    1052    1071
0    1179    7    2    5    1100    1152    1116    1089    1134
0    1181    7    1    2    1089    1111
0    1182    7    1    3    1100    1089    1128
0    1183    7    1    4    1116    1089    1145    1100
0    1184    7    1    5    1134    1116    1089    1160    1100
0    1188    7    1    2    1100    1128
0    1189    7    1    3    1116    1145    1100
0    1190    7    1    4    1134    1116    1160    1100
0    1191    7    1    5    4    1152    1116    1134    1100
0    1192    7    1    2    1145    1116
0    1193    7    1    3    1134    1116    1160
0    1194    7    1    4    4    1152    1116    1134
0    1195    7    1    2    1134    1160
0    1196    7    1    3    4    1152    1134
0    1197    7    1    2    4    1152
0    1437    7    2    4    1422    1307    1289    1278
0    1442    7    1    2    1289    1318
0    1443    7    1    3    1307    1324    1289
0    1444    7    1    3    1422    1307    1289
0    1445    7    1    2    1289    1318
0    1446    7    1    3    1307    1324    1289
0    1447    7    1    2    1307    1324
0    1451    7    2    5    1430    1390    1365    1344    1332
0    1454    7    1    2    1332    1359
0    1455    7    1    3    1344    1332    1382
0    1456    7    1    4    1365    1332    1404    1344
0    1457    7    1    5    1390    1365    1332    1412    1344
0    1465    7    1    2    1344    1382
0    1466    7    1    3    1365    1404    1344
0    1467    7    1    4    1390    1365    1412    1344
0    1468    7    1    4    1430    1365    1344    1390
0    1469    7    1    2    1344    1382
0    1470    7    1    3    1365    1404    1344
0    1471    7    1    4    1390    1365    1412    1344
0    1472    7    1    2    1365    1404
0    1473    7    1    3    1390    1365    1412
0    1474    7    1    3    1430    1365    1390
0    1475    7    1    2    1365    1404
0    1476    7    1    3    1390    1365    1412
0    1477    7    1    2    1390    1412
0    1481    7    1    2    1422    1307
0    1482    7    1    2    1430    1390
0    1764    5    1    1    1758
0    1843    7    2    4    1712    1758    1730    1704
0    1850    7    1    3    1730    1749    1712
0    1851    7    1    3    1758    1730    1712
0    1853    7    1    3    1749    1730    1712
0    1854    7    1    2    1730    1749
0    1855    7    1    2    1758    1730
0    1856    7    1    2    1730    1749
0    1857    7    2    5    1778    1829    1794    1767    1812
0    1859    7    1    2    1767    1789
0    1860    7    1    3    1778    1767    1806
0    1861    7    1    4    1794    1767    1823    1778
0    1862    7    1    5    1812    1794    1767    1837    1778
0    1867    7    1    3    1794    1823    1778
0    1868    7    1    4    1812    1794    1837    1778
0    1869    7    1    5    54    1829    1794    1812    1778
0    1870    7    1    2    1823    1794
0    1871    7    1    3    1812    1794    1837
0    1872    7    1    4    54    1829    1794    1812
0    1873    7    1    2    1812    1837
0    1874    7    1    3    54    1829    1812
0    1878    6    2    2    1876    1877
0    2113    7    2    4    2099    1984    1966    1958
0    2120    7    1    3    1984    2001    1966
0    2121    7    1    3    2099    1984    1966
0    2123    7    1    3    1984    2001    1966
0    2124    7    1    2    1984    2001
0    2128    7    2    5    2106    2067    2042    2021    2009
0    2131    7    1    2    2009    2036
0    2132    7    1    3    2021    2009    2059
0    2133    7    1    4    2042    2009    2081    2021
0    2134    7    1    5    2067    2042    2009    2089    2021
0    2143    7    1    3    2042    2081    2021
0    2144    7    1    4    2067    2042    2089    2021
0    2145    7    1    4    2106    2042    2021    2067
0    2147    7    1    3    2042    2081    2021
0    2148    7    1    4    2067    2042    2089    2021
0    2149    7    1    2    2042    2081
0    2150    7    1    3    2067    2042    2089
0    2151    7    1    3    2106    2042    2067
0    2152    7    1    2    2042    2081
0    2153    7    1    3    2067    2042    2089
0    2154    7    1    2    2067    2089
0    2158    7    1    2    2099    1984
0    2159    7    1    2    2106    2067
0    3449    5    2    1    3445
0    3458    5    2    1    3454
0    3472    5    2    1    3468
0    3481    5    2    1    3477
2    3497    1    3463
2    3501    1    3463
2    3505    1    3486
2    3509    1    3486
0    3531    6    1    2    5239    5242
0    5428    5    1    1    5422
0    3967    6    1    2    5422    5429
2    4191    1    1152
2    4199    1    1023
2    4207    1    1023
2    4215    1    1034
2    4223    1    1034
2    4231    1    1052
2    4239    1    1052
2    4247    1    1089
2    4255    1    1100
2    4263    1    1116
2    4271    1    1134
2    4371    1    1422
2    4381    1    1307
2    4391    1    1278
2    4401    1    1289
2    4429    1    1422
2    4439    1    1307
2    4449    1    1278
2    4459    1    1289
2    4497    1    1430
2    4507    1    1390
2    4517    1    1332
2    4527    1    1365
2    4537    1    1344
2    4547    1    1344
2    4585    1    1430
2    4595    1    1390
2    4605    1    1332
2    4615    1    1365
2    4719    1    1730
2    4727    1    1730
2    4735    1    1767
2    4751    1    1794
2    4759    1    1812
2    4835    1    2099
2    4845    1    1984
2    4893    1    2099
2    4903    1    1984
2    4961    1    2067
2    4971    1    2009
2    4981    1    2042
2    5049    1    2067
2    5059    1    2009
2    5069    1    2042
0    5222    5    1    1    5216
0    5223    5    1    1    5219
0    5232    5    1    1    5226
0    5233    5    1    1    5229
0    5294    6    1    2    5289    5292
0    5395    6    1    2    5386    5393
0    589    3    1    4    1286    1439    1440    1441
0    616    3    1    4    3167    1845    1846    1847
0    619    3    1    4    1031    1168    1169    1170
0    627    3    1    4    3167    2115    2116    2117
0    1185    3    2    5    1097    1181    1182    1183    1184
0    1448    3    2    2    1318    1447
0    1458    3    3    5    1341    1454    1455    1456    1457
0    1478    3    2    2    1404    1477
0    1863    3    2    5    1775    1859    1860    1861    1862
0    4747    5    1    1    4743
0    2125    3    2    2    1995    2124
0    2135    3    3    5    2018    2131    2132    2133    2134
0    2155    3    2    2    2081    2154
0    4995    5    1    1    4991
0    5005    5    1    1    5001
0    3533    6    2    2    3531    3532
0    3921    5    1    1    3918
0    3925    5    1    1    3922
0    3929    5    1    1    3926
0    3933    5    1    1    3930
0    3943    7    1    3    3862    3853    3918
0    3946    7    1    3    3866    3857    3922
0    3949    7    1    3    3883    3874    3926
0    3952    7    1    3    3887    3878    3930
0    3966    6    1    2    5425    5428
0    4107    6    2    2    4104    132
0    4196    3    2    4    1046    1171    1172    1173
0    4204    4    2    3    1046    1174    1175
0    4212    3    2    3    1064    1176    1177
0    4220    4    2    2    1064    1178
0    4244    3    2    5    1111    1188    1189    1190    1191
0    4252    3    2    4    1128    1192    1193    1194
0    4260    3    2    3    1145    1195    1196
0    4268    3    2    2    1160    1197
0    4361    3    2    4    1301    1442    1443    1444
0    4419    4    2    3    1301    1445    1446
0    4467    3    2    4    1382    1472    1473    1474
0    4487    3    2    5    1359    1465    1466    1467    1468
0    4555    4    2    3    1382    1475    1476
0    4575    4    2    4    1359    1469    1470    1471
0    4684    3    2    4    1724    1849    1850    1851
0    4692    4    2    3    1724    1852    1853
0    4700    3    2    3    1742    1854    1855
0    4708    4    2    2    1742    1856
0    4732    3    2    5    1789    1866    1867    1868    1869
0    4740    3    2    4    1806    1870    1871    1872
0    4748    3    2    3    1823    1873    1874
0    4825    3    2    4    1978    2119    2120    2121
0    4883    4    2    3    1978    2122    2123
0    4928    3    2    4    2059    2149    2150    2151
0    4941    3    2    5    2036    2142    2143    2144    2145
0    5009    4    2    3    2059    2152    2153
0    5029    4    2    4    2036    2146    2147    2148
0    5224    6    1    2    5219    5222
0    5225    6    1    2    5216    5223
0    5234    6    1    2    5229    5232
0    5235    6    1    2    5226    5233
0    5376    6    2    2    5294    5295
0    5417    6    2    2    5394    5395
0    576    5    1    1    1878
3    588    7    0    2    1437    1451
3    615    7    0    2    1843    1857
3    626    7    0    2    2113    2128
3    632    7    0    2    1166    1179
0    1198    6    1    2    4191    4194
0    4195    5    1    1    4191
0    4203    5    1    1    4199
0    4211    5    1    1    4207
0    4219    5    1    1    4215
0    4227    5    1    1    4223
0    1217    6    1    2    4231    4234
0    4235    5    1    1    4231
0    1221    6    1    2    4239    4242
0    4243    5    1    1    4239
0    1224    7    1    2    1179    4
0    4251    5    1    1    4247
0    4259    5    1    1    4255
0    4267    5    1    1    4263
0    4275    5    1    1    4271
0    1453    5    1    1    1451
0    4405    5    1    1    4401
0    4463    5    1    1    4459
0    4541    5    1    1    4537
0    4551    5    1    1    4547
0    1895    6    1    2    4719    4722
0    4723    5    1    1    4719
0    1899    6    1    2    4727    4730
0    4731    5    1    1    4727
0    1902    7    1    2    1857    54
0    4739    5    1    1    4735
0    4755    5    1    1    4751
0    1929    6    1    2    4759    4762
0    4763    5    1    1    4759
0    2130    5    1    1    2128
0    3500    5    1    1    3497
0    3504    5    1    1    3501
0    3508    5    1    1    3505
0    3512    5    1    1    3509
0    3520    7    1    3    3454    3445    3497
0    3523    7    1    3    3458    3449    3501
0    3526    7    1    3    3477    3468    3505
0    3529    7    1    3    3481    3472    3509
3    1002    1    0    1    3533
0    3837    7    1    3    1878    3795    3823
0    3942    7    1    3    3857    3862    3921
0    3945    7    1    3    3853    3866    3925
0    3948    7    1    3    3878    3883    3929
0    3951    7    1    3    3874    3887    3933
0    3968    6    2    2    3966    3967
0    4375    5    1    1    4371
0    4385    5    1    1    4381
0    4395    5    1    1    4391
0    4433    5    1    1    4429
0    4443    5    1    1    4439
0    4453    5    1    1    4449
0    4501    5    1    1    4497
0    4511    5    1    1    4507
0    4521    5    1    1    4517
0    4531    5    1    1    4527
0    4619    5    1    1    4615
0    4589    5    1    1    4585
0    4599    5    1    1    4595
0    4609    5    1    1    4605
0    4839    5    1    1    4835
0    4849    5    1    1    4845
0    4897    5    1    1    4893
0    4907    5    1    1    4903
0    4965    5    1    1    4961
0    4975    5    1    1    4971
0    4985    5    1    1    4981
0    5073    5    1    1    5069
0    5053    5    1    1    5049
0    5063    5    1    1    5059
0    5247    6    2    2    5224    5225
0    5255    6    2    2    5234    5235
0    590    7    1    2    1437    1458
0    617    7    1    2    1863    1843
0    620    7    1    2    1185    1166
0    628    7    1    2    2113    2135
0    3535    5    1    1    3533
0    1199    6    1    2    4188    4195
0    4202    5    1    1    4196
0    1204    6    1    2    4196    4203
0    4210    5    1    1    4204
0    1207    6    1    2    4204    4211
0    4218    5    1    1    4212
0    1211    6    1    2    4212    4219
0    4226    5    1    1    4220
0    1214    6    1    2    4220    4227
0    1218    6    1    2    4228    4235
0    1222    6    1    2    4236    4243
0    1225    3    5    2    1185    1224
0    4250    5    1    1    4244
0    1237    6    1    2    4244    4251
0    4258    5    1    1    4252
0    1242    6    1    2    4252    4259
0    4266    5    1    1    4260
0    1247    6    1    2    4260    4267
0    4274    5    1    1    4268
0    1252    6    1    2    4268    4275
0    1462    5    2    1    1458
0    4690    5    1    1    4684
0    1882    6    1    2    4684    4691
0    4698    5    1    1    4692
0    1885    6    1    2    4692    4699
0    4706    5    1    1    4700
0    1889    6    1    2    4700    4707
0    4714    5    1    1    4708
0    1892    6    1    2    4708    4715
0    1896    6    1    2    4716    4723
0    1900    6    1    2    4724    4731
0    1903    3    5    2    1863    1902
0    4738    5    1    1    4732
0    1915    6    1    2    4732    4739
0    4746    5    1    1    4740
0    1920    6    1    2    4740    4747
0    4754    5    1    1    4748
0    1925    6    1    2    4748    4755
0    1930    6    1    2    4756    4763
0    2139    5    2    1    2135
0    3519    7    1    3    3449    3454    3500
0    3522    7    1    3    3445    3458    3504
0    3525    7    1    3    3472    3477    3508
0    3528    7    1    3    3468    3481    3512
0    3848    3    5    3    3836    3837    3838
0    3944    4    1    2    3942    3943
0    3947    4    1    2    3945    3946
0    3950    4    1    2    3948    3949
0    3953    4    1    2    3951    3952
0    5421    5    1    1    5417
3    1004    1    0    1    3968
0    4111    7    1    2    4104    4107
0    4112    7    1    2    4107    132
0    4351    3    2    2    1448    1481
0    4365    5    1    1    4361
0    4409    5    2    1    1448
0    4423    5    1    1    4419
0    4471    5    1    1    4467
0    4472    6    1    2    4467    4470
0    4477    3    2    2    1478    1482
0    4491    5    1    1    4487
0    4559    5    1    1    4555
0    4560    6    1    2    4555    4558
0    4565    5    2    1    1478
0    4579    5    1    1    4575
0    4815    3    2    2    2125    2158
0    4829    5    1    1    4825
0    4873    5    2    1    2125
0    4887    5    1    1    4883
0    4931    3    2    2    2155    2159
0    4934    5    1    1    4928
0    4945    5    1    1    4941
0    5013    5    1    1    5009
0    5014    6    1    2    5009    5012
0    5019    5    2    1    2155
0    5033    5    1    1    5029
0    5382    5    1    1    5376
0    5385    6    1    2    5376    5383
3    591    3    0    2    589    590
3    618    3    0    2    616    617
3    621    3    0    2    619    620
3    629    3    0    2    627    628
0    3970    5    1    1    3968
0    1200    6    2    2    1198    1199
0    1203    6    1    2    4199    4202
0    1206    6    1    2    4207    4210
0    1210    6    1    2    4215    4218
0    1213    6    1    2    4223    4226
0    1219    6    1    2    1217    1218
0    1223    6    1    2    1221    1222
0    1236    6    1    2    4247    4250
0    1241    6    1    2    4255    4258
0    1246    6    1    2    4263    4266
0    1251    6    1    2    4271    4274
0    1881    6    1    2    4687    4690
0    1884    6    1    2    4695    4698
0    1888    6    1    2    4703    4706
0    1891    6    1    2    4711    4714
0    1897    6    1    2    1895    1896
0    1901    6    1    2    1899    1900
0    1914    6    1    2    4735    4738
0    1919    6    1    2    4743    4746
0    1924    6    1    2    4751    4754
0    1931    6    2    2    1929    1930
0    3521    4    1    2    3519    3520
0    3524    4    1    2    3522    3523
0    3527    4    1    2    3525    3526
0    3530    4    1    2    3528    3529
0    5251    5    1    1    5247
0    5259    5    1    1    5255
0    4113    3    3    2    4111    4112
0    4473    6    1    2    4464    4471
0    4561    6    1    2    4552    4559
0    5015    6    1    2    5006    5013
0    5384    6    1    2    5379    5382
0    5406    6    2    2    3947    3944
0    5414    6    2    2    3953    3950
0    1664    7    1    3    3848    1621    1645
0    2335    7    1    3    3848    2293    2316
0    718    7    1    3    3848    2430    2454
3    822    5    0    1    3848
0    855    7    1    3    3848    2488    2512
0    1205    6    1    2    1203    1204
0    1208    6    1    2    1206    1207
0    1212    6    1    2    1210    1211
0    1215    6    1    2    1213    1214
0    1220    5    1    1    1219
0    1231    5    4    1    1225
0    1238    6    2    2    1236    1237
0    1243    6    2    2    1241    1242
0    1248    6    2    2    1246    1247
0    1253    6    2    2    1251    1252
0    1272    7    1    2    1225    1086
0    1483    7    2    2    1462    1453
0    1883    6    1    2    1881    1882
0    1886    6    1    2    1884    1885
0    1890    6    1    2    1888    1889
0    1893    6    1    2    1891    1892
0    1898    5    1    1    1897
0    1909    5    4    1    1903
0    1916    6    2    2    1914    1915
0    1921    6    2    2    1919    1920
0    1926    6    2    2    1924    1925
0    1953    7    1    2    1903    1764
0    2160    7    2    2    2139    2130
0    4355    5    1    1    4351
0    4356    6    1    2    4351    4354
0    4413    5    1    1    4409
0    4414    6    1    2    4409    4412
0    4474    6    2    2    4472    4473
0    4481    5    1    1    4477
0    4562    6    2    2    4560    4561
0    4569    5    1    1    4565
0    4819    5    1    1    4815
0    4820    6    1    2    4815    4818
0    4877    5    1    1    4873
0    4878    6    1    2    4873    4876
0    4935    5    1    1    4931
0    4936    6    1    2    4931    4934
0    5016    6    2    2    5014    5015
0    5023    5    1    1    5019
0    5244    6    2    2    3524    3521
0    5252    6    2    2    3530    3527
0    5409    6    2    2    5384    5385
0    566    5    1    1    1200
0    577    5    1    1    1931
0    3733    7    1    3    4113    3724    3721
0    1209    5    1    1    1208
0    1216    5    1    1    1215
0    1257    7    1    2    1225    1205
0    1262    7    1    2    1225    1212
0    1267    7    1    2    1225    1220
0    1887    5    1    1    1886
0    1894    5    1    1    1893
0    1935    7    1    2    1903    1883
0    1943    7    1    2    1903    1890
0    1948    7    1    2    1903    1898
0    3779    7    1    3    1200    3737    3765
0    3840    7    1    3    1931    3795    3823
0    5412    5    1    1    5406
0    5420    5    1    1    5414
0    3964    6    1    2    5414    5421
0    4357    6    1    2    4348    4355
0    4415    6    1    2    4406    4413
0    4821    6    1    2    4812    4819
0    4879    6    1    2    4870    4877
0    4937    6    1    2    4928    4935
0    567    5    1    1    1253
0    568    5    1    1    1248
0    569    5    1    1    1243
0    570    5    1    1    1238
0    578    5    1    1    1926
0    579    5    1    1    1921
0    580    5    1    1    1916
0    1256    7    1    2    1209    1231
0    1261    7    1    2    1216    1231
0    1266    7    1    2    1223    1231
0    1271    7    1    2    1080    1231
0    1486    5    1    1    1483
0    1934    7    1    2    1887    1909
0    1942    7    1    2    1894    1909
0    1947    7    1    2    1901    1909
0    1952    7    1    2    1758    1909
0    2163    5    1    1    2160
0    5250    5    1    1    5244
0    3537    6    1    2    5244    5251
0    5258    5    1    1    5252
0    3542    6    1    2    5252    5259
0    3782    7    1    3    1253    3737    3765
0    3785    7    1    3    1248    3737    3765
0    3788    7    1    3    1243    3737    3765
0    3790    3    5    3    3778    3779    3780
0    3843    7    1    3    1926    3795    3823
0    3846    7    1    3    1921    3795    3823
0    3849    3    5    3    3839    3840    3841
0    3960    6    1    2    5409    5412
0    5413    5    1    1    5409
0    3963    6    1    2    5417    5420
0    4010    7    1    3    1238    3972    3998
0    4068    7    1    3    1916    4030    4056
0    4358    6    2    2    4356    4357
0    4416    6    2    2    4414    4415
0    4480    5    1    1    4474
0    4483    6    1    2    4474    4481
0    4568    5    1    1    4562
0    4571    6    1    2    4562    4569
0    4822    6    2    2    4820    4821
0    4880    6    2    2    4878    4879
0    4938    6    2    2    4936    4937
0    5022    5    1    1    5016
0    5025    6    1    2    5016    5023
0    1258    3    2    2    1256    1257
0    1263    3    2    2    1261    1262
0    1268    3    2    2    1266    1267
0    1273    3    2    2    1271    1272
0    1936    3    6    2    1934    1935
0    1944    3    2    2    1942    1943
0    1949    3    2    2    1947    1948
0    1954    3    2    2    1952    1953
0    3536    6    1    2    5247    5250
0    3541    6    1    2    5255    5258
0    3791    3    5    3    3781    3782    3783
0    3792    3    5    3    3784    3785    3786
0    3793    3    5    3    3787    3788    3789
0    3850    3    5    3    3842    3843    3844
0    3851    3    5    3    3845    3846    3847
0    3961    6    1    2    5406    5413
0    3965    6    2    2    3963    3964
0    4024    3    5    3    4009    4010    4011
0    4082    3    5    3    4067    4068    4069
0    4482    6    1    2    4477    4480
0    4570    6    1    2    4565    4568
0    5024    6    1    2    5019    5022
0    1666    7    1    3    3790    1609    1645
0    1670    7    1    3    3849    1621    1645
0    2337    7    1    3    3790    2281    2316
0    2341    7    1    3    3849    2293    2316
0    719    7    1    3    3790    2418    2454
0    758    7    1    3    3849    2430    2454
0    798    7    1    3    3849    2488    2512
3    838    5    0    1    3849
0    856    7    1    3    3790    2476    2512
3    861    5    0    1    3790
0    3538    6    2    2    3536    3537
0    3543    6    2    2    3541    3542
0    3962    6    2    2    3960    3961
0    4364    5    1    1    4358
0    4367    6    1    2    4358    4365
0    4422    5    1    1    4416
0    4425    6    1    2    4416    4423
0    4484    6    2    2    4482    4483
0    4572    6    2    2    4570    4571
0    4828    5    1    1    4822
0    4831    6    1    2    4822    4829
0    4886    5    1    1    4880
0    4889    6    1    2    4880    4887
0    4944    5    1    1    4938
0    4947    6    1    2    4938    4945
0    5026    6    2    2    5024    5025
0    571    5    1    1    1273
0    572    5    1    1    1268
0    573    5    1    1    1263
0    574    5    1    1    1258
0    581    5    1    1    1954
0    582    5    1    1    1949
0    583    5    1    1    1944
0    584    5    1    1    1936
3    623    5    0    1    1936
0    1576    7    1    3    4082    1540    1564
0    1578    7    1    3    4024    1528    1564
0    659    3    1    4    1664    1666    1667    1668
0    1672    7    1    3    3791    1609    1645
0    1676    7    1    3    3850    1621    1645
0    1678    7    1    3    3792    1609    1645
0    1682    7    1    3    3851    1621    1645
0    1684    7    1    3    3793    1609    1645
0    2250    7    1    3    4082    2215    2238
0    2252    7    1    3    4024    2203    2238
0    691    3    1    4    2335    2337    2338    2339
0    2343    7    1    3    3791    2281    2316
0    2347    7    1    3    3850    2293    2316
0    2349    7    1    3    3792    2281    2316
0    2353    7    1    3    3851    2293    2316
0    2355    7    1    3    3793    2281    2316
3    722    3    0    4    718    719    720    721
0    743    7    1    3    4082    3570    3594
0    744    7    1    3    4024    3558    3594
0    748    7    1    3    3851    2430    2454
0    749    7    1    3    3793    2418    2454
0    753    7    1    3    3850    2430    2454
0    754    7    1    3    3792    2418    2454
0    759    7    1    3    3791    2418    2454
0    783    7    1    3    4082    3672    3696
0    784    7    1    3    4024    3660    3696
0    788    7    1    3    3851    2488    2512
0    789    7    1    3    3793    2476    2512
0    793    7    1    3    3850    2488    2512
0    794    7    1    3    3792    2476    2512
0    799    7    1    3    3791    2476    2512
0    3735    7    1    3    1936    3724    3717
3    832    5    0    1    4082
3    834    5    0    1    3851
3    836    5    0    1    3850
0    3835    5    1    1    3965
3    859    3    0    4    855    856    857    858
3    871    5    0    1    4024
3    873    5    0    1    3793
3    875    5    0    1    3792
3    877    5    0    1    3791
3    998    1    0    1    3538
3    1000    1    0    1    3543
0    3651    7    1    2    3965    3632
0    4013    7    1    3    1273    3972    3998
0    4016    7    1    3    1268    3972    3998
0    4019    7    1    3    1263    3972    3998
0    4022    7    1    3    1258    3972    3998
0    4071    7    1    3    1954    4030    4056
0    4074    7    1    3    1949    4030    4056
0    4077    7    1    3    1944    4030    4056
0    4080    7    1    3    1936    4030    4056
0    4096    6    2    2    4113    1936
0    4366    6    1    2    4361    4364
0    4424    6    1    2    4419    4422
0    4830    6    1    2    4825    4828
0    4888    6    1    2    4883    4886
0    4946    6    1    2    4941    4944
3    575    7    0    9    566    567    568    569    570    571    572    573    574
3    585    7    0    9    576    577    578    579    580    581    582    583    584
0    640    3    1    4    1576    1578    1579    1580
3    661    7    0    2    659    1606
0    662    3    1    4    1670    1672    1673    1674
0    665    3    1    4    1676    1678    1679    1680
0    668    3    1    4    1682    1684    1685    1686
0    674    3    1    4    2250    2252    2253    2254
3    693    7    0    2    691    2279
0    694    3    1    4    2341    2343    2344    2345
0    697    3    1    4    2347    2349    2350    2351
0    700    3    1    4    2353    2355    2356    2357
3    747    3    0    4    743    744    745    746
3    752    3    0    4    748    749    750    751
3    757    3    0    4    753    754    755    756
3    762    3    0    4    758    759    760    761
3    787    3    0    4    783    784    785    786
3    792    3    0    4    788    789    790    791
3    797    3    0    4    793    794    795    796
3    802    3    0    4    798    799    800    801
0    817    3    1    4    3731    3733    3734    3735
0    839    7    1    3    3835    3803    3823
0    3540    5    1    1    3538
0    3545    5    1    1    3543
0    3777    5    1    1    3962
0    3648    7    1    2    3962    3632
0    4025    3    5    3    4012    4013    4014
0    4026    3    5    3    4015    4016    4017
0    4027    3    5    3    4018    4019    4020
0    4028    3    5    3    4021    4022    4023
0    4083    3    5    3    4070    4071    4072
0    4084    3    5    3    4073    4074    4075
0    4085    3    5    3    4076    4077    4078
0    4086    3    5    3    4079    4080    4081
0    4368    6    2    2    4366    4367
0    4426    6    2    2    4424    4425
0    4490    5    1    1    4484
0    4493    6    1    2    4484    4491
0    4578    5    1    1    4572
0    4581    6    1    2    4572    4579
0    4832    6    2    2    4830    4831
0    4890    6    2    2    4888    4889
0    4948    6    2    2    4946    4947
0    5032    5    1    1    5026
0    5035    6    1    2    5026    5033
3    642    7    0    2    640    1526
3    664    7    0    2    662    1606
3    667    7    0    2    665    1606
3    670    7    0    2    668    1606
3    676    7    0    2    674    2202
3    696    7    0    2    694    2279
3    699    7    0    2    697    2279
3    702    7    0    2    700    2279
0    811    7    1    2    4113    4096
0    812    7    1    2    4096    1936
3    818    7    0    2    816    817
0    853    7    1    5    562    3540    3545    3535    3970
0    878    7    1    3    3777    3745    3765
0    4492    6    1    2    4487    4490
0    4580    6    1    2    4575    4578
0    5034    6    1    2    5029    5032
0    1582    7    1    3    4083    1540    1564
0    1584    7    1    3    4025    1528    1564
0    1588    7    1    3    4084    1540    1564
0    1590    7    1    3    4026    1528    1564
0    1594    7    1    3    4085    1540    1564
0    1596    7    1    3    4027    1528    1564
0    1600    7    1    3    4086    1540    1564
0    1602    7    1    3    4028    1528    1564
0    2256    7    1    3    4083    2215    2238
0    2258    7    1    3    4025    2203    2238
0    2262    7    1    3    4084    2215    2238
0    2264    7    1    3    4026    2203    2238
0    2268    7    1    3    4085    2215    2238
0    2270    7    1    3    4027    2203    2238
0    2274    7    1    3    4086    2215    2238
0    2276    7    1    3    4028    2203    2238
0    708    7    1    3    4086    3672    3696
0    709    7    1    3    4028    3660    3696
0    723    7    1    3    4086    3570    3594
0    724    7    1    3    4028    3558    3594
0    728    7    1    3    4085    3570    3594
0    729    7    1    3    4027    3558    3594
0    733    7    1    3    4084    3570    3594
0    734    7    1    3    4026    3558    3594
0    738    7    1    3    4083    3570    3594
0    739    7    1    3    4025    3558    3594
0    768    7    1    3    4085    3672    3696
0    769    7    1    3    4027    3660    3696
0    773    7    1    3    4084    3672    3696
0    774    7    1    3    4026    3660    3696
0    778    7    1    3    4083    3672    3696
0    779    7    1    3    4025    3660    3696
3    813    3    0    2    811    812
3    824    5    0    1    4086
3    826    5    0    1    4085
3    828    5    0    1    4084
3    830    5    0    1    4083
3    854    7    0    3    852    853    245
3    863    5    0    1    4028
3    865    5    0    1    4027
3    867    5    0    1    4026
3    869    5    0    1    4025
0    4374    5    1    1    4368
0    4377    6    1    2    4368    4375
0    4432    5    1    1    4426
0    4435    6    1    2    4426    4433
0    4494    6    2    2    4492    4493
0    4582    6    2    2    4580    4581
0    4838    5    1    1    4832
0    4841    6    1    2    4832    4839
0    4896    5    1    1    4890
0    4899    6    1    2    4890    4897
0    4954    5    1    1    4948
0    4957    6    1    2    4948    4955
0    5036    6    2    2    5034    5035
0    643    3    1    4    1582    1584    1585    1586
0    646    3    1    4    1588    1590    1591    1592
0    649    3    1    4    1594    1596    1597    1598
0    652    3    1    4    1600    1602    1603    1604
0    677    3    1    4    2256    2258    2259    2260
0    680    3    1    4    2262    2264    2265    2266
0    683    3    1    4    2268    2270    2271    2272
0    686    3    1    4    2274    2276    2277    2278
3    712    3    0    4    708    709    710    711
3    727    3    0    4    723    724    725    726
3    732    3    0    4    728    729    730    731
3    737    3    0    4    733    734    735    736
3    742    3    0    4    738    739    740    741
3    772    3    0    4    768    769    770    771
3    777    3    0    4    773    774    775    776
3    782    3    0    4    778    779    780    781
0    4376    6    1    2    4371    4374
0    4434    6    1    2    4429    4432
0    4840    6    1    2    4835    4838
0    4898    6    1    2    4893    4896
0    4956    6    1    2    4951    4954
3    645    7    0    2    643    1526
3    648    7    0    2    646    1526
3    651    7    0    2    649    1526
3    654    7    0    2    652    1526
3    679    7    0    2    677    2202
3    682    7    0    2    680    2202
3    685    7    0    2    683    2202
3    688    7    0    2    686    2202
0    4378    6    2    2    4376    4377
0    4436    6    2    2    4434    4435
0    4500    5    1    1    4494
0    4503    6    1    2    4494    4501
0    4588    5    1    1    4582
0    4591    6    1    2    4582    4589
0    4842    6    2    2    4840    4841
0    4900    6    2    2    4898    4899
0    4958    6    2    2    4956    4957
0    5042    5    1    1    5036
0    5045    6    1    2    5036    5043
0    4502    6    1    2    4497    4500
0    4590    6    1    2    4585    4588
0    5044    6    1    2    5039    5042
0    4384    5    1    1    4378
0    4387    6    1    2    4378    4385
0    4442    5    1    1    4436
0    4445    6    1    2    4436    4443
0    4504    6    2    2    4502    4503
0    4592    6    2    2    4590    4591
0    4848    5    1    1    4842
0    4851    6    1    2    4842    4849
0    4906    5    1    1    4900
0    4909    6    1    2    4900    4907
0    4964    5    1    1    4958
0    4967    6    1    2    4958    4965
0    5046    6    2    2    5044    5045
0    4386    6    1    2    4381    4384
0    4444    6    1    2    4439    4442
0    4850    6    1    2    4845    4848
0    4908    6    1    2    4903    4906
0    4966    6    1    2    4961    4964
0    4388    6    2    2    4386    4387
0    4446    6    2    2    4444    4445
0    4510    5    1    1    4504
0    4513    6    1    2    4504    4511
0    4598    5    1    1    4592
0    4601    6    1    2    4592    4599
0    4852    6    2    2    4850    4851
0    4910    6    2    2    4908    4909
0    4968    6    2    2    4966    4967
0    5052    5    1    1    5046
0    5055    6    1    2    5046    5053
0    4512    6    1    2    4507    4510
0    4600    6    1    2    4595    4598
0    5054    6    1    2    5049    5052
0    4394    5    1    1    4388
0    4397    6    1    2    4388    4395
0    4452    5    1    1    4446
0    4455    6    1    2    4446    4453
0    4514    6    2    2    4512    4513
0    4602    6    2    2    4600    4601
0    4858    5    1    1    4852
0    4861    6    1    2    4852    4859
0    4916    5    1    1    4910
0    4919    6    1    2    4910    4917
0    4974    5    1    1    4968
0    4977    6    1    2    4968    4975
0    5056    6    2    2    5054    5055
0    4396    6    1    2    4391    4394
0    4454    6    1    2    4449    4452
0    4860    6    1    2    4855    4858
0    4918    6    1    2    4913    4916
0    4976    6    1    2    4971    4974
0    4398    6    2    2    4396    4397
0    4456    6    2    2    4454    4455
0    4520    5    1    1    4514
0    4523    6    1    2    4514    4521
0    4608    5    1    1    4602
0    4611    6    1    2    4602    4609
0    4862    6    2    2    4860    4861
0    4920    6    2    2    4918    4919
0    4978    6    2    2    4976    4977
0    5062    5    1    1    5056
0    5065    6    1    2    5056    5063
0    4522    6    1    2    4517    4520
0    4610    6    1    2    4605    4608
0    5064    6    1    2    5059    5062
0    4404    5    1    1    4398
0    1488    6    1    2    4398    4405
0    4462    5    1    1    4456
0    1493    6    1    2    4456    4463
0    4868    5    1    1    4862
0    2165    6    1    2    4862    4869
0    4926    5    1    1    4920
0    2170    6    1    2    4920    4927
0    4524    6    2    2    4522    4523
0    4612    6    2    2    4610    4611
0    4984    5    1    1    4978
0    4987    6    1    2    4978    4985
0    5066    6    2    2    5064    5065
0    1487    6    1    2    4401    4404
0    1492    6    1    2    4459    4462
0    2164    6    1    2    4865    4868
0    2169    6    1    2    4923    4926
0    4986    6    1    2    4981    4984
0    1489    6    2    2    1487    1488
0    1494    6    2    2    1492    1493
0    2166    6    2    2    2164    2165
0    2171    6    2    2    2169    2170
0    4530    5    1    1    4524
0    4533    6    1    2    4524    4531
0    4618    5    1    1    4612
0    4543    6    1    2    4612    4619
0    4988    6    2    2    4986    4987
0    5072    5    1    1    5066
0    4997    6    1    2    5066    5073
0    4532    6    1    2    4527    4530
0    4542    6    1    2    4615    4618
0    4996    6    1    2    5069    5072
0    1513    7    1    3    1494    1462    1502
0    1514    7    1    3    1489    1458    1502
0    1515    7    1    3    1494    1483    1497
0    1516    7    1    3    1489    1486    1497
0    4994    5    1    1    4988
0    2184    6    1    2    4988    4995
0    2190    7    1    3    2171    2139    2179
0    2191    7    1    3    2166    2135    2179
0    2192    7    1    3    2171    2160    2174
0    2193    7    1    3    2166    2163    2174
0    4534    6    2    2    4532    4533
0    4544    6    2    2    4542    4543
0    4998    6    2    2    4996    4997
0    2183    6    1    2    4991    4994
0    4620    3    2    4    1513    1514    1515    1516
0    5074    3    2    4    2190    2191    2192    2193
0    4540    5    1    1    4534
0    1507    6    1    2    4534    4541
0    4550    5    1    1    4544
0    1510    6    1    2    4544    4551
0    2185    6    1    2    2183    2184
0    5004    5    1    1    4998
0    2187    6    1    2    4998    5005
0    1506    6    1    2    4537    4540
0    1509    6    1    2    4547    4550
0    4626    5    1    1    4620
0    2186    6    1    2    5001    5004
0    2195    7    1    2    2174    2185
0    5080    5    1    1    5074
0    1508    6    1    2    1506    1507
0    1511    6    1    2    1509    1510
0    2188    6    1    2    2186    2187
0    1512    5    1    1    1511
0    1518    7    1    2    1497    1508
0    2189    5    1    1    2188
0    1517    7    1    2    1512    1502
0    2194    7    1    2    2189    2179
0    4623    3    2    2    1517    1518
0    5077    3    2    2    2194    2195
0    1519    6    1    2    4623    4626
0    4627    5    1    1    4623
0    2196    6    1    2    5077    5080
0    5081    5    1    1    5077
0    1520    6    1    2    4620    4627
0    2197    6    1    2    5074    5081
0    1521    6    2    2    1519    1520
0    2198    6    2    2    2196    2197
0    840    7    1    3    2198    3795    3823
0    879    7    1    3    1521    3737    3765
0    1524    5    1    1    1521
0    2201    5    1    1    2198
3    843    3    0    4    839    840    841    842
3    882    3    0    4    878    879    880    881
0    3649    7    1    2    1524    3628
0    3652    7    1    2    2201    3628
0    3657    3    2    2    3648    3649
0    3658    3    2    2    3651    3652
0    3636    7    1    2    3657    3622
0    3639    7    1    2    3658    3622
0    3642    7    1    2    3657    3622
0    3645    7    1    2    3658    3622
0    3653    3    2    2    3636    3637
0    3654    3    2    2    3639    3640
0    3655    3    2    2    3642    3643
0    3656    3    2    2    3645    3646
0    763    7    1    3    3656    2430    2454
0    764    7    1    3    3655    2418    2454
0    803    7    1    3    3656    2488    2512
0    804    7    1    3    3655    2476    2512
0    1657    7    1    3    3654    1621    1645
0    1659    7    1    3    3653    1609    1645
0    2328    7    1    3    3654    2293    2316
0    2330    7    1    3    3653    2281    2316
0    1662    3    1    4    1657    1659    1660    1661
0    2333    3    1    4    2328    2330    2331    2332
3    767    3    0    4    763    764    765    766
3    807    3    0    4    803    804    805    806
0    657    7    1    2    1662    1606
0    689    7    1    2    2333    2279
3    658    5    0    1    657
3    690    5    0    1    689
