1 1 0 1 0
1 2 0 1 0
1 3 0 2 0
1 4 0 2 0
1 5 0 2 0
1 6 0 2 0
2 7 1 3
2 8 1 4
2 9 1 5
2 10 1 6
0 11 7 1 2 1 2
0 12 2 1 2 3 4
0 13 2 1 2 5 6
0 14 8 1 2 7 8
0 15 8 1 2 9 10
0 16 2 1 2 12 13
0 17 8 1 2 14 15
0 18 2 1 2 11 16
3 19 2 1 2 18 17