1    153    0    1    0
1    1459    0    1    0
1    188    0    1    0
1    165    0    1    0
1    191    0    1    0
1    44    0    1    0
1    3705    0    1    0
1    4400    0    1    0
1    157    0    1    0
1    74    0    1    0
1    228    0    1    0
1    234    0    1    0
1    3717    0    1    0
1    216    0    1    0
1    109    0    1    0
1    3698    0    1    0
1    85    0    1    0
1    12    0    1    0
1    230    0    1    0
1    88    0    1    0
1    1486    0    1    0
1    156    0    1    0
1    118    0    1    0
1    223    0    1    0
1    64    0    1    0
1    163    0    1    0
1    187    0    1    0
1    4528    0    1    0
1    184    0    1    0
1    2247    0    1    0
1    213    0    1    0
1    2208    0    1    0
1    75    0    1    0
1    164    0    1    0
1    214    0    1    0
1    203    0    1    0
1    181    0    1    0
1    221    0    1    0
1    226    0    1    0
1    240    0    1    0
1    81    0    1    0
1    207    0    1    0
1    205    0    1    0
1    219    0    1    0
1    38    0    1    0
1    26    0    1    0
1    3749    0    1    0
1    112    0    1    0
1    167    0    1    0
1    151    0    1    0
1    1496    0    1    0
1    171    0    1    0
1    50    0    1    0
1    235    0    1    0
1    172    0    1    0
1    2204    0    1    0
1    1    0    1    0
1    1197    0    1    0
1    23    0    1    0
1    160    0    1    0
1    4405    0    1    0
1    56    0    1    0
1    62    0    1    0
1    154    0    1    0
1    222    0    1    0
1    3723    0    1    0
1    3743    0    1    0
1    3729    0    1    0
1    138    0    1    0
1    158    0    1    0
1    183    0    1    0
1    232    0    1    0
1    35    0    1    0
1    77    0    1    0
1    87    0    1    0
1    113    0    1    0
1    173    0    1    0
1    180    0    1    0
1    176    0    1    0
1    70    0    1    0
1    4526    0    1    0
1    57    0    1    0
1    103    0    1    0
1    59    0    1    0
1    86    0    1    0
1    195    0    1    0
1    141    0    1    0
1    80    0    1    0
1    94    0    1    0
1    1469    0    1    0
1    4437    0    1    0
1    159    0    1    0
1    218    0    1    0
1    2253    0    1    0
1    166    0    1    0
1    9    0    1    0
1    134    0    1    0
1    63    0    1    0
1    197    0    1    0
1    206    0    1    0
1    100    0    1    0
1    124    0    1    0
1    127    0    1    0
1    54    0    1    0
1    15    0    1    0
1    220    0    1    0
1    196    0    1    0
1    76    0    1    0
1    84    0    1    0
1    192    0    1    0
1    41    0    1    0
1    237    0    1    0
1    1462    0    1    0
1    4394    0    1    0
1    2211    0    1    0
1    73    0    1    0
1    152    0    1    0
1    97    0    1    0
1    175    0    1    0
1    4427    0    1    0
1    2236    0    1    0
1    4432    0    1    0
1    233    0    1    0
1    135    0    1    0
1    190    0    1    0
1    202    0    1    0
1    66    0    1    0
1    2239    0    1    0
1    4410    0    1    0
1    182    0    1    0
1    225    0    1    0
1    79    0    1    0
1    147    0    1    0
1    61    0    1    0
1    168    0    1    0
1    177    0    1    0
1    2230    0    1    0
1    53    0    1    0
1    60    0    1    0
1    5    0    1    0
1    47    0    1    0
1    2256    0    1    0
1    199    0    1    0
1    58    0    1    0
1    83    0    1    0
1    215    0    1    0
1    2218    0    1    0
1    1480    0    1    0
1    229    0    1    0
1    161    0    1    0
1    4420    0    1    0
1    3737    0    1    0
1    115    0    1    0
1    55    0    1    0
1    4393    0    1    0
1    212    0    1    0
1    339    0    1    0
1    201    0    1    0
1    231    0    1    0
1    29    0    1    0
1    114    0    1    0
1    179    0    1    0
1    186    0    1    0
1    198    0    1    0
1    69    0    1    0
1    193    0    1    0
1    3711    0    1    0
1    209    0    1    0
1    1455    0    1    0
1    162    0    1    0
1    150    0    1    0
1    4415    0    1    0
1    208    0    1    0
1    82    0    1    0
1    236    0    1    0
1    170    0    1    0
1    18    0    1    0
1    110    0    1    0
1    106    0    1    0
1    204    0    1    0
1    178    0    1    0
1    238    0    1    0
1    130    0    1    0
1    89    0    1    0
1    239    0    1    0
1    3701    0    1    0
1    32    0    1    0
1    1492    0    1    0
1    200    0    1    0
1    174    0    1    0
1    224    0    1    0
1    227    0    1    0
1    189    0    1    0
1    144    0    1    0
1    111    0    1    0
1    194    0    1    0
1    185    0    1    0
1    78    0    1    0
1    211    0    1    0
1    210    0    1    0
1    155    0    1    0
1    133    0    1    0
1    121    0    1    0
1    2224    0    1    0
1    65    0    1    0
1    169    0    1    0
1    217    0    1    0
3    2    1    0    1    1
3    3    1    0    1    1
0    400    5    1    1    57
0    1184    7    2    2    134    133
3    450    1    0    1    1459
3    448    1    0    1    1469
3    444    1    0    1    1480
3    442    1    0    1    1486
3    440    1    0    1    1492
3    438    1    0    1    1496
0    1501    7    2    4    162    172    188    199
3    496    1    0    1    2208
3    494    1    0    1    2218
3    492    1    0    1    2224
3    490    1    0    1    2230
3    488    1    0    1    2236
3    486    1    0    1    2239
3    484    1    0    1    2247
3    482    1    0    1    2253
3    480    1    0    1    2256
0    2857    7    2    4    150    184    228    240
3    560    1    0    1    3698
3    542    1    0    1    3701
3    558    1    0    1    3705
3    556    1    0    1    3711
3    554    1    0    1    3717
3    552    1    0    1    3723
3    550    1    0    1    3729
3    548    1    0    1    3737
3    546    1    0    1    3743
3    544    1    0    1    3749
3    540    1    0    1    4393
3    538    1    0    1    4400
3    536    1    0    1    4405
3    534    1    0    1    4410
3    532    1    0    1    4415
3    530    1    0    1    4420
3    528    1    0    1    4427
3    526    1    0    1    4432
3    524    1    0    1    4437
0    4442    7    2    4    183    182    185    186
0    4514    7    2    4    210    152    218    230
3    279    5    0    1    15
0    401    5    1    1    5
2    573    1    1
0    574    5    2    1    5
0    575    5    2    1    5
0    1178    5    4    1    2236
0    1186    5    4    1    2253
0    1192    5    4    1    2256
2    1198    1    38
2    1205    1    15
0    1206    6    3    2    12    9
0    1207    6    3    2    12    9
2    1210    1    38
0    1458    5    1    1    1455
0    1461    5    1    1    1459
3    436    1    0    1    1462
0    1464    5    6    1    1462
0    1471    5    5    1    1469
2    1475    1    106
0    1482    5    5    1    1480
0    1488    5    5    1    1486
0    1495    5    1    1    1492
0    1499    5    1    1    1496
0    1500    5    1    1    106
2    1503    1    18
2    1512    1    18
0    1518    7    1    2    4528    1492
2    1524    1    18
0    1535    5    4    1    18
0    1541    6    4    2    4528    1496
0    2207    5    1    1    2204
0    2210    5    1    1    2208
3    478    1    0    1    2211
0    2213    5    6    1    2211
0    2220    5    5    1    2218
0    2226    5    5    1    2224
0    2232    5    5    1    2230
0    2238    5    1    1    2236
0    2241    5    7    1    2239
0    2249    5    5    1    2247
0    2255    5    1    1    2253
0    2258    5    1    1    2256
2    2828    1    4526
0    3700    5    1    1    3698
0    3703    5    2    1    3701
0    3707    5    5    1    3705
0    3713    5    5    1    3711
0    3719    5    5    1    3717
0    3725    5    5    1    3723
0    3731    5    7    1    3729
0    3739    5    5    1    3737
0    3745    5    5    1    3743
0    3751    5    5    1    3749
0    4121    5    1    1    4393
3    522    1    0    1    4394
0    4396    5    6    1    4394
0    4402    5    5    1    4400
0    4407    5    5    1    4405
0    4412    5    5    1    4410
0    4417    5    5    1    4415
0    4422    5    7    1    4420
0    4429    5    5    1    4427
0    4434    5    5    1    4432
0    4439    5    5    1    4437
2    4833    1    4526
3    402    6    0    2    400    401
3    404    5    0    1    2857
3    406    5    0    1    4514
3    408    5    0    1    4442
3    410    5    0    1    1501
0    2876    7    1    2    2857    4514
0    2878    7    1    2    4442    1501
3    432    1    0    1    573
3    446    1    0    1    1475
0    1519    5    6    1    1518
0    2871    7    1    2    4528    1458
0    2883    6    2    2    4528    2207
0    280    7    1    2    1184    575
3    284    6    0    2    1197    574
3    286    5    0    1    1205
3    289    6    0    2    1197    574
3    292    6    0    2    1184    575
3    341    5    0    1    1205
0    4839    5    1    1    4833
2    572    1    573
2    581    1    1206
2    587    1    1512
2    601    1    1206
2    606    1    1512
2    650    1    1206
2    657    1    1512
2    671    1    1207
2    678    1    1503
0    777    7    4    2    1541    1198
0    1115    7    1    2    1541    1198
2    1336    1    1512
2    1350    1    1503
0    1477    5    4    1    1475
0    1507    5    4    1    1503
0    1514    5    2    1    1512
0    1530    5    4    1    1524
2    2259    1    1535
0    2833    5    3    1    2828
0    2872    5    2    1    2871
2    2886    1    1207
2    2892    1    1503
2    2905    1    1207
2    2909    1    1503
2    3622    1    1524
2    3635    1    1524
2    3755    1    1535
2    4640    1    1524
2    4653    1    1524
2    4873    1    1541
2    4876    1    1198
2    4881    1    1488
2    4889    1    1482
2    4905    1    1471
2    4916    1    1198
2    4921    1    1464
2    5175    1    1541
2    5178    1    1198
2    5186    1    1198
2    5191    1    1488
2    5199    1    1482
2    5215    1    1471
2    5223    1    1464
2    5393    1    1192
2    5401    1    1186
2    5409    1    2249
2    5417    1    1178
2    5425    1    2232
2    5433    1    2226
2    5441    1    2220
2    5449    1    2241
2    5457    1    2213
2    5745    1    1192
2    5753    1    1186
2    5761    1    2249
2    5769    1    2241
2    5777    1    1178
2    5785    1    2232
2    5793    1    2226
2    5801    1    2220
2    5809    1    2213
2    5865    1    3751
2    5873    1    3745
2    5881    1    3739
2    5889    1    3731
2    5897    1    3725
2    5905    1    3719
2    5913    1    3713
2    5921    1    3707
2    5985    1    3751
2    5993    1    3745
2    6001    1    3739
2    6009    1    3725
2    6017    1    3719
2    6025    1    3713
2    6033    1    3707
2    6041    1    3731
2    6514    1    1210
2    6554    1    1210
2    6567    1    4439
2    6575    1    4434
2    6583    1    4429
2    6591    1    4422
2    6599    1    4417
2    6607    1    4412
2    6615    1    4407
2    6623    1    4402
2    6631    1    4396
2    6853    1    4439
2    6861    1    4434
2    6869    1    4429
2    6877    1    4417
2    6885    1    4412
2    6893    1    4407
2    6901    1    4402
2    6909    1    4422
2    6917    1    4396
3    281    5    0    1    280
3    453    1    0    1    572
0    784    7    5    2    1519    1198
0    1014    7    2    2    1198    1519
0    3221    7    1    2    2883    1210
2    4913    1    1519
0    4929    4    2    2    1519    1198
2    5183    1    1519
0    5231    4    2    2    1198    1519
2    6511    1    2883
3    278    7    0    2    163    572
0    615    7    1    2    170    587
0    594    5    5    1    587
0    611    5    3    1    606
0    617    7    1    2    169    587
0    619    7    1    2    168    587
0    621    7    1    2    167    587
0    623    7    1    2    166    606
0    625    7    1    2    165    606
0    627    7    1    2    164    606
0    664    5    5    1    657
0    685    5    5    1    678
0    691    7    1    2    177    657
0    693    7    1    2    176    657
0    695    7    1    2    175    657
0    697    7    1    2    174    657
0    699    7    1    2    173    657
0    701    7    1    2    157    678
0    703    7    1    2    156    678
0    705    7    1    2    155    678
0    707    7    1    2    154    678
0    709    7    1    2    153    678
0    4879    5    1    1    4873
0    4880    5    1    1    4876
0    4887    5    1    1    4881
0    4895    5    1    1    4889
0    4911    5    1    1    4905
0    4920    5    1    1    4916
0    4927    5    1    1    4921
0    5181    5    1    1    5175
0    5182    5    1    1    5178
0    5190    5    1    1    5186
0    5197    5    1    1    5191
0    5205    5    1    1    5199
0    5221    5    1    1    5215
0    5229    5    1    1    5223
0    1343    5    5    1    1336
0    1357    5    5    1    1350
0    1364    7    1    2    181    1336
0    1366    7    1    2    171    1336
0    1368    7    1    2    180    1336
0    1370    7    1    2    179    1336
0    1372    7    1    2    178    1336
0    1374    7    1    2    161    1350
0    1376    7    1    2    151    1350
0    1378    7    1    2    160    1350
0    1380    7    1    2    159    1350
0    1382    7    1    2    158    1350
0    5399    5    1    1    5393
0    5407    5    1    1    5401
0    5415    5    1    1    5409
0    5423    5    1    1    5417
0    5431    5    1    1    5425
0    5439    5    1    1    5433
0    5447    5    1    1    5441
0    5455    5    1    1    5449
0    5463    5    1    1    5457
0    5751    5    1    1    5745
0    5759    5    1    1    5753
0    5767    5    1    1    5761
0    5775    5    1    1    5769
0    5783    5    1    1    5777
0    5791    5    1    1    5785
0    5799    5    1    1    5793
0    5807    5    1    1    5801
0    5815    5    1    1    5809
2    2019    1    1514
2    2032    1    1507
2    2117    1    1514
2    2130    1    1507
0    2266    5    5    1    2259
2    2272    1    1507
0    2286    7    1    2    44    2259
0    2288    7    1    2    41    2259
0    2290    7    1    2    29    2259
0    2292    7    1    2    26    2259
0    2294    7    1    2    23    2259
0    5871    5    1    1    5865
0    5879    5    1    1    5873
0    5887    5    1    1    5881
0    5895    5    1    1    5889
0    5903    5    1    1    5897
0    5911    5    1    1    5905
0    5919    5    1    1    5913
0    5927    5    1    1    5921
0    5991    5    1    1    5985
0    5999    5    1    1    5993
0    6007    5    1    1    6001
0    6015    5    1    1    6009
0    6023    5    1    1    6017
0    6031    5    1    1    6025
0    6039    5    1    1    6033
0    6047    5    1    1    6041
0    2899    5    5    1    2892
0    2914    5    3    1    2909
0    2919    7    1    2    209    2892
0    2921    7    1    2    216    2892
0    2923    7    1    2    215    2892
0    2925    7    1    2    214    2892
0    2927    7    1    2    213    2909
0    2929    7    1    2    212    2909
0    2931    7    1    2    211    2909
0    6518    5    1    1    6514
0    3173    7    1    2    2872    1210
0    6558    5    1    1    6554
0    6573    5    1    1    6567
0    6581    5    1    1    6575
0    6589    5    1    1    6583
0    6597    5    1    1    6591
0    6605    5    1    1    6599
0    6613    5    1    1    6607
0    6621    5    1    1    6615
0    6629    5    1    1    6623
0    6637    5    1    1    6631
0    3629    5    5    1    3622
0    3642    5    5    1    3635
0    3649    7    1    2    1461    3622
0    3651    7    1    2    1464    3622
0    3653    7    1    2    1471    3622
0    3655    7    1    2    1500    3622
0    3657    7    1    2    1482    3622
0    3659    7    1    2    1488    3635
0    3661    7    1    2    1495    3635
0    3663    7    1    2    1499    3635
0    3762    5    5    1    3755
2    3768    1    1507
0    3782    7    1    2    47    3755
0    3784    7    1    2    35    3755
0    3786    7    1    2    32    3755
0    3788    7    1    2    50    3755
0    3790    7    1    2    66    3755
0    6859    5    1    1    6853
0    6867    5    1    1    6861
0    6875    5    1    1    6869
0    6883    5    1    1    6877
0    6891    5    1    1    6885
0    6899    5    1    1    6893
0    6907    5    1    1    6901
0    6915    5    1    1    6909
0    6923    5    1    1    6917
2    4094    1    1530
2    4107    1    1530
2    4444    1    1530
2    4457    1    1530
0    4647    5    5    1    4640
0    4660    5    5    1    4653
0    4667    7    1    2    2210    4640
0    4669    7    1    2    2213    4640
0    4671    7    1    2    2220    4640
0    4673    7    1    2    2226    4640
0    4675    7    1    2    2232    4640
0    4677    7    1    2    2238    4653
0    4679    7    1    2    2241    4653
0    4681    7    1    2    2249    4653
0    4683    7    1    2    2255    4653
0    4685    7    1    2    2258    4653
2    4897    1    1477
2    5207    1    1477
2    6551    1    2872
0    763    6    1    2    4876    4879
0    764    6    1    2    4873    4880
0    4919    5    1    1    4913
0    886    6    1    2    4913    4920
0    1005    6    1    2    5178    5181
0    1006    6    1    2    5175    5182
0    5189    5    1    1    5183
0    1018    6    1    2    5183    5190
0    5237    5    1    1    5231
0    6517    5    1    1    6511
0    3169    6    1    2    6511    6518
0    4935    5    1    1    4929
2    4970    1    784
2    5239    1    1014
0    577    3    1    2    594    615
0    616    3    1    2    594    587
0    618    3    1    2    594    617
0    620    3    1    2    594    619
0    622    3    1    2    594    621
0    624    3    1    2    611    623
0    626    3    1    2    611    625
0    628    3    1    2    611    627
0    692    3    1    2    664    691
0    694    3    1    2    664    693
0    696    3    1    2    664    695
0    698    3    1    2    664    697
0    700    3    1    2    664    699
0    702    3    1    2    685    701
0    704    3    1    2    685    703
0    706    3    1    2    685    705
0    708    3    1    2    685    707
0    710    3    1    2    685    709
0    765    6    9    2    763    764
0    4903    5    1    1    4897
0    885    6    1    2    4916    4919
0    1007    6    4    2    1005    1006
0    1017    6    1    2    5186    5189
0    5213    5    1    1    5207
0    1363    7    1    2    141    1343
0    1365    7    1    2    147    1343
0    1367    7    1    2    138    1343
0    1369    7    1    2    144    1343
0    1371    7    1    2    135    1343
0    1373    7    1    2    141    1357
0    1375    7    1    2    147    1357
0    1377    7    1    2    138    1357
0    1379    7    1    2    144    1357
0    1381    7    1    2    135    1357
0    2026    5    5    1    2019
0    2039    5    5    1    2032
0    2046    7    1    2    103    2019
0    2048    7    1    2    130    2019
0    2050    7    1    2    127    2019
0    2052    7    1    2    124    2019
0    2054    7    1    2    100    2019
0    2056    7    1    2    103    2032
0    2058    7    1    2    130    2032
0    2060    7    1    2    127    2032
0    2062    7    1    2    124    2032
0    2064    7    1    2    100    2032
0    2124    5    5    1    2117
0    2137    5    5    1    2130
0    2144    7    1    2    115    2117
0    2146    7    1    2    118    2117
0    2148    7    1    2    97    2117
0    2150    7    1    2    94    2117
0    2152    7    1    2    121    2117
0    2154    7    1    2    115    2130
0    2156    7    1    2    118    2130
0    2158    7    1    2    97    2130
0    2160    7    1    2    94    2130
0    2162    7    1    2    121    2130
0    2279    5    5    1    2272
0    2285    7    1    2    208    2266
0    2287    7    1    2    198    2266
0    2289    7    1    2    207    2266
0    2291    7    1    2    206    2266
0    2293    7    1    2    205    2266
0    2296    7    1    2    44    2272
0    2298    7    1    2    41    2272
0    2300    7    1    2    29    2272
0    2302    7    1    2    26    2272
0    2304    7    1    2    23    2272
0    2918    3    1    2    2899    2892
0    2920    3    1    2    2899    2919
0    2922    3    1    2    2899    2921
0    2924    3    1    2    2899    2923
0    2926    3    1    2    2899    2925
0    2928    3    1    2    2914    2927
0    2930    3    1    2    2914    2929
0    2932    3    1    2    2914    2931
0    3168    6    1    2    6514    6517
0    6557    5    1    1    6551
0    3211    6    1    2    6551    6558
0    3648    7    1    2    114    3629
0    3650    7    1    2    113    3629
0    3652    7    1    2    111    3629
0    3654    7    1    2    87    3629
0    3656    7    1    2    112    3629
0    3658    7    1    2    88    3642
0    3660    7    1    2    1455    3642
0    3662    7    1    2    2204    3642
0    3665    7    1    2    3703    3642
0    3666    7    1    2    70    3642
0    3775    5    5    1    3768
0    3781    7    1    2    193    3762
0    3783    7    1    2    192    3762
0    3785    7    1    2    191    3762
0    3787    7    1    2    190    3762
0    3789    7    1    2    189    3762
0    3792    7    1    2    47    3768
0    3794    7    1    2    35    3768
0    3796    7    1    2    32    3768
0    3798    7    1    2    50    3768
0    3800    7    1    2    66    3768
0    4101    5    5    1    4094
0    4114    5    5    1    4107
0    4123    7    1    2    58    4094
0    4126    7    1    2    77    4094
0    4129    7    1    2    78    4094
0    4132    7    1    2    59    4094
0    4135    7    1    2    81    4094
0    4138    7    1    2    80    4107
0    4141    7    1    2    79    4107
0    4144    7    1    2    60    4107
0    4147    7    1    2    61    4107
0    4150    7    1    2    62    4107
0    4451    5    5    1    4444
0    4464    5    5    1    4457
0    4471    7    1    2    69    4444
0    4473    7    1    2    70    4444
0    4475    7    1    2    74    4444
0    4477    7    1    2    76    4444
0    4479    7    1    2    75    4444
0    4481    7    1    2    73    4457
0    4483    7    1    2    53    4457
0    4485    7    1    2    54    4457
0    4487    7    1    2    55    4457
0    4489    7    1    2    56    4457
0    4666    7    1    2    82    4647
0    4668    7    1    2    65    4647
0    4670    7    1    2    83    4647
0    4672    7    1    2    84    4647
0    4674    7    1    2    85    4647
0    4676    7    1    2    64    4660
0    4678    7    1    2    63    4660
0    4680    7    1    2    86    4660
0    4682    7    1    2    109    4660
0    4684    7    1    2    110    4660
0    579    7    1    2    577    581
0    629    7    3    2    616    581
0    633    7    3    2    618    581
0    637    7    3    2    620    581
0    641    7    3    2    622    581
0    645    7    3    2    624    601
0    711    7    3    2    692    650
0    715    7    3    2    694    650
0    719    7    3    2    696    650
0    723    7    3    2    698    650
0    727    7    3    2    700    650
0    731    7    5    2    702    671
0    737    7    7    2    704    671
0    745    7    5    2    706    671
0    751    7    5    2    708    671
0    757    7    5    2    710    671
0    887    6    5    2    885    886
0    1019    6    3    2    1017    1018
0    5245    5    1    1    5239
0    1383    3    3    2    1365    1366
0    1387    3    3    2    1367    1368
0    1391    3    3    2    1369    1370
0    1395    3    3    2    1371    1372
0    1399    3    6    2    1375    1376
0    1406    3    5    2    1377    1378
0    1412    3    5    2    1379    1380
0    1418    3    5    2    1381    1382
0    2305    3    2    2    2287    2288
0    2308    3    3    2    2289    2290
0    2312    3    3    2    2291    2292
0    2316    3    3    2    2293    2294
0    2933    7    6    2    2920    2886
0    2938    7    5    2    2922    2886
0    2942    7    5    2    2924    2886
0    2946    7    5    2    2926    2886
0    2950    7    5    2    2928    2905
0    3170    6    2    2    3168    3169
0    3210    6    1    2    6554    6557
0    3667    3    3    2    3650    3651
0    3670    3    3    2    3652    3653
0    3673    3    3    2    3654    3655
0    3676    3    3    2    3656    3657
0    3679    3    3    2    3658    3659
0    3682    3    5    2    3665    3635
0    3686    3    2    2    3666    3635
0    3801    3    3    2    3781    3782
0    3804    3    3    2    3783    3784
0    3807    3    3    2    3785    3786
0    3810    3    3    2    3787    3788
0    3813    3    3    2    3789    3790
0    4525    7    1    2    2918    2886
0    4686    3    3    2    4668    4669
0    4689    3    3    2    4670    4671
0    4692    3    3    2    4672    4673
0    4695    3    3    2    4674    4675
0    4698    3    3    2    4676    4677
0    4701    3    3    2    4678    4679
0    4704    3    3    2    4680    4681
0    4707    3    3    2    4682    4683
0    4710    3    3    2    4684    4685
0    4976    5    1    1    4970
0    5271    7    2    2    2932    2905
0    5274    7    2    2    2930    2905
0    5305    7    2    2    628    601
0    5308    7    2    2    626    601
0    5318    3    2    2    1373    1374
0    6690    3    2    2    3648    3649
0    6711    3    2    2    3662    3663
0    6714    3    2    2    3660    3661
0    7252    3    2    2    2285    2286
0    7296    3    2    2    1363    1364
0    7466    3    2    2    4666    4667
0    907    7    1    2    765    784
0    913    7    1    2    765    784
0    915    7    1    2    765    784
0    916    7    1    2    765    784
0    1116    7    1    2    1007    1014
0    2045    7    1    2    204    2026
0    2047    7    1    2    203    2026
0    2049    7    1    2    202    2026
0    2051    7    1    2    201    2026
0    2053    7    1    2    200    2026
0    2055    7    1    2    235    2039
0    2057    7    1    2    234    2039
0    2059    7    1    2    233    2039
0    2061    7    1    2    232    2039
0    2063    7    1    2    231    2039
0    2143    7    1    2    197    2124
0    2145    7    1    2    187    2124
0    2147    7    1    2    196    2124
0    2149    7    1    2    195    2124
0    2151    7    1    2    194    2124
0    2153    7    1    2    227    2137
0    2155    7    1    2    217    2137
0    2157    7    1    2    226    2137
0    2159    7    1    2    225    2137
0    2161    7    1    2    224    2137
0    2295    7    1    2    239    2279
0    2297    7    1    2    229    2279
0    2299    7    1    2    238    2279
0    2301    7    1    2    237    2279
0    2303    7    1    2    236    2279
0    3212    6    1    2    3210    3211
0    3791    7    1    2    223    3775
0    3793    7    1    2    222    3775
0    3795    7    1    2    221    3775
0    3797    7    1    2    220    3775
0    3799    7    1    2    219    3775
0    4122    7    1    2    4121    4101
0    4125    7    1    2    4396    4101
0    4128    7    1    2    4402    4101
0    4131    7    1    2    4407    4101
0    4134    7    1    2    4412    4101
0    4137    7    1    2    4417    4114
0    4140    7    1    2    4422    4114
0    4143    7    1    2    4429    4114
0    4146    7    1    2    4434    4114
0    4149    7    1    2    4439    4114
0    4470    7    1    2    3700    4451
0    4472    7    1    2    3703    4451
0    4474    7    1    2    3707    4451
0    4476    7    1    2    3713    4451
0    4478    7    1    2    3719    4451
0    4480    7    1    2    3725    4464
0    4482    7    1    2    3731    4464
0    4484    7    1    2    3739    4464
0    4486    7    1    2    3745    4464
0    4488    7    1    2    3751    4464
2    4962    1    765
2    5003    1    765
2    5234    1    1007
2    5242    1    1007
0    5250    5    2    1    4525
0    5284    5    2    1    579
0    802    7    1    2    1488    2950
0    821    7    3    2    1482    2946
0    845    7    5    2    1477    2942
0    868    7    6    2    1471    2938
0    877    7    7    2    1464    2933
0    902    7    3    2    887    765
0    908    3    3    2    777    907
0    914    7    1    2    887    765
0    917    3    2    2    777    916
0    953    7    1    2    887    765
0    1023    5    1    1    1019
0    1035    7    1    2    1488    2950
0    1050    7    2    2    1482    2946
0    1068    7    3    2    1477    2942
0    1086    7    4    2    1471    2938
0    1102    7    5    2    1464    2933
0    1108    7    3    2    1019    1007
0    1117    3    3    2    1115    1116
0    5322    5    1    1    5318
0    1553    7    1    2    1192    757
0    1567    7    3    2    1186    751
0    1584    7    4    2    2249    745
0    1590    7    5    2    2241    737
0    1606    7    1    2    1178    731
0    1624    7    3    2    2232    1418
0    1647    7    5    2    2226    1412
0    1669    7    6    2    2220    1406
0    1677    7    7    2    2213    1399
0    1802    7    1    2    1192    757
0    1816    7    3    2    1186    751
0    1834    7    5    2    2249    745
0    1841    7    6    2    737    2241
0    1866    7    1    2    1178    731
0    1880    7    2    2    2232    1418
0    1897    7    3    2    2226    1412
0    1914    7    4    2    2220    1406
0    1929    7    5    2    2213    1399
0    2065    3    3    2    2045    2046
0    2069    3    3    2    2047    2048
0    2073    3    3    2    2049    2050
0    2077    3    3    2    2051    2052
0    2081    3    3    2    2053    2054
0    2085    3    5    2    2055    2056
0    2091    3    7    2    2057    2058
0    2099    3    5    2    2059    2060
0    2105    3    5    2    2061    2062
0    2111    3    5    2    2063    2064
0    2163    3    3    2    2145    2146
0    2167    3    3    2    2147    2148
0    2171    3    3    2    2149    2150
0    2175    3    3    2    2151    2152
0    2179    3    6    2    2155    2156
0    2186    3    5    2    2157    2158
0    2192    3    5    2    2159    2160
0    2198    3    5    2    2161    2162
0    2320    3    2    2    2297    2298
0    2323    3    5    2    2299    2300
0    2329    3    5    2    2301    2302
0    2335    3    5    2    2303    2304
0    2962    7    1    2    4710    727
0    2970    7    1    2    4707    723
0    2977    7    1    2    4704    719
0    2979    7    1    2    4701    715
0    2989    7    1    2    4698    711
0    2998    7    1    2    4695    1395
0    3006    7    1    2    4692    1391
0    3013    7    1    2    4689    1387
0    3015    7    1    2    4686    1383
0    3183    7    1    2    3679    645
0    3192    7    1    2    3676    641
0    3200    7    1    2    3673    637
0    3207    7    1    2    3670    633
0    3209    7    1    2    3667    629
0    3216    7    3    2    3212    3170
0    3222    7    1    2    3170    3173
0    6694    5    1    1    6690
0    3695    7    2    2    1535    2305
0    3816    3    5    2    3791    3792
0    3821    3    7    2    3793    3794
0    3828    3    5    2    3795    3796
0    3833    3    5    2    3797    3798
0    3838    3    5    2    3799    3800
0    4151    3    3    2    4125    4126
0    4154    3    3    2    4128    4129
0    4157    3    3    2    4131    4132
0    4160    3    3    2    4134    4135
0    4163    3    3    2    4137    4138
0    4166    3    3    2    4140    4141
0    4169    3    3    2    4143    4144
0    4172    3    3    2    4146    4147
0    4175    3    3    2    4149    4150
0    7256    5    1    1    7252
0    7300    5    1    1    7296
0    4490    3    3    2    4474    4475
0    4493    3    3    2    4476    4477
0    4496    3    3    2    4478    4479
0    4499    3    3    2    4480    4481
0    4502    3    3    2    4482    4483
0    4505    3    3    2    4484    4485
0    4508    3    3    2    4486    4487
0    4511    3    3    2    4488    4489
0    7470    5    1    1    7466
2    4884    1    2950
2    4892    1    2946
2    4900    1    2942
2    4908    1    2938
2    4924    1    2933
2    4952    1    887
0    4983    4    2    2    777    915
2    4993    1    887
0    5011    4    2    2    1464    2933
2    5194    1    2950
2    5202    1    2946
2    5210    1    2942
2    5218    1    2938
2    5226    1    2933
2    5247    1    2933
2    5255    1    2942
2    5258    1    2938
2    5263    1    2950
2    5266    1    2946
0    5277    5    1    1    5271
0    5278    5    1    1    5274
2    5281    1    629
2    5289    1    637
2    5292    1    633
2    5297    1    645
2    5300    1    641
0    5311    5    1    1    5305
0    5312    5    1    1    5308
2    5315    1    1399
2    5323    1    1412
2    5326    1    1406
2    5331    1    731
2    5334    1    1418
2    5339    1    745
2    5342    1    737
2    5349    1    757
2    5352    1    751
2    5396    1    757
2    5404    1    751
2    5412    1    745
2    5420    1    731
2    5428    1    1418
2    5436    1    1412
2    5444    1    1406
2    5452    1    737
2    5460    1    1399
0    5465    4    2    2    2241    737
0    5581    4    2    2    2213    1399
2    5748    1    757
2    5756    1    751
2    5764    1    745
2    5772    1    737
2    5780    1    731
2    5788    1    1418
2    5796    1    1412
2    5804    1    1406
2    5812    1    1399
0    5849    4    2    2    737    2241
2    5929    1    3682
2    6049    1    3682
2    6367    1    4710
2    6370    1    727
2    6375    1    4707
2    6378    1    723
2    6383    1    4704
2    6386    1    719
2    6391    1    4698
2    6394    1    711
2    6399    1    4695
2    6402    1    1395
2    6407    1    4692
2    6410    1    1391
2    6415    1    4689
2    6418    1    1387
2    6423    1    4701
2    6426    1    715
2    6431    1    4686
2    6434    1    1383
2    6442    1    3813
2    6450    1    3810
2    6458    1    3807
2    6466    1    3801
2    6498    1    3804
2    6519    1    3679
2    6522    1    645
2    6527    1    3676
2    6530    1    641
2    6535    1    3673
2    6538    1    637
2    6543    1    3670
2    6546    1    633
2    6559    1    3667
2    6562    1    629
2    6687    1    3667
2    6695    1    3673
2    6698    1    3670
2    6703    1    3679
2    6706    1    3676
0    6717    5    1    1    6711
0    6718    5    1    1    6714
0    6724    3    2    2    2153    2154
0    6768    3    2    2    2295    2296
0    7208    3    2    2    2143    2144
2    7221    1    3801
2    7229    1    3807
2    7232    1    3804
2    7239    1    3813
2    7242    1    3810
2    7249    1    2305
2    7257    1    2312
2    7260    1    2308
2    7268    1    2316
2    7293    1    1383
2    7301    1    1391
2    7304    1    1387
2    7309    1    711
2    7312    1    1395
2    7317    1    719
2    7320    1    715
2    7327    1    727
2    7330    1    723
2    7396    1    2316
2    7404    1    2312
2    7412    1    2308
2    7425    1    3686
2    7463    1    4686
2    7471    1    4692
2    7474    1    4689
2    7479    1    4698
2    7482    1    4695
2    7487    1    4704
2    7490    1    4701
2    7497    1    4710
2    7500    1    4707
0    7507    3    2    2    4472    4473
0    7510    3    2    2    4470    4471
0    7554    3    2    2    4122    4123
0    1152    6    1    2    5234    5237
0    5238    5    1    1    5234
0    1156    6    1    2    5242    5245
0    5246    5    1    1    5242
0    5254    5    1    1    5250
0    5288    5    1    1    5284
0    3223    3    3    2    3221    3222
0    4942    3    2    3    777    913    914
0    4966    5    1    1    4962
0    5007    5    1    1    5003
0    5279    6    1    2    5274    5277
0    5280    6    1    2    5271    5278
0    5313    6    1    2    5308    5311
0    5314    6    1    2    5305    5312
0    6719    6    1    2    6714    6717
0    6720    6    1    2    6711    6718
0    790    6    1    2    4884    4887
0    4888    5    1    1    4884
0    803    6    1    2    4892    4895
0    4896    5    1    1    4892
0    825    6    1    2    4900    4903
0    4904    5    1    1    4900
0    851    6    1    2    4908    4911
0    4912    5    1    1    4908
0    893    6    1    2    4924    4927
0    4928    5    1    1    4924
0    906    5    1    1    902
0    912    5    1    1    908
0    1024    6    1    2    5194    5197
0    5198    5    1    1    5194
0    1036    6    1    2    5202    5205
0    5206    5    1    1    5202
0    1053    6    1    2    5210    5213
0    5214    5    1    1    5210
0    1072    6    1    2    5218    5221
0    5222    5    1    1    5218
0    1091    6    1    2    5226    5229
0    5230    5    1    1    5226
0    1112    5    1    1    1108
0    1121    5    1    1    1117
0    1153    6    1    2    5231    5238
0    1157    6    1    2    5239    5246
0    5253    5    1    1    5247
0    1216    6    1    2    5247    5254
0    5261    5    1    1    5255
0    5262    5    1    1    5258
0    5269    5    1    1    5263
0    5270    5    1    1    5266
0    5287    5    1    1    5281
0    1239    6    1    2    5281    5288
0    5295    5    1    1    5289
0    5296    5    1    1    5292
0    5303    5    1    1    5297
0    5304    5    1    1    5300
0    5321    5    1    1    5315
0    1262    6    1    2    5315    5322
0    5329    5    1    1    5323
0    5330    5    1    1    5326
0    5337    5    1    1    5331
0    5338    5    1    1    5334
0    1544    6    1    2    5396    5399
0    5400    5    1    1    5396
0    1554    6    1    2    5404    5407
0    5408    5    1    1    5404
0    1571    6    1    2    5412    5415
0    5416    5    1    1    5412
0    1596    6    1    2    5420    5423
0    5424    5    1    1    5420
0    1607    6    1    2    5428    5431
0    5432    5    1    1    5428
0    1628    6    1    2    5436    5439
0    5440    5    1    1    5436
0    1653    6    1    2    5444    5447
0    5448    5    1    1    5444
0    1685    6    1    2    5452    5455
0    5456    5    1    1    5452
0    1693    6    1    2    5460    5463
0    5464    5    1    1    5460
0    1793    6    1    2    5748    5751
0    5752    5    1    1    5748
0    1803    6    1    2    5756    5759
0    5760    5    1    1    5756
0    1820    6    1    2    5764    5767
0    5768    5    1    1    5764
0    1848    6    1    2    5772    5775
0    5776    5    1    1    5772
0    1857    6    1    2    5780    5783
0    5784    5    1    1    5780
0    1867    6    1    2    5788    5791
0    5792    5    1    1    5788
0    1883    6    1    2    5796    5799
0    5800    5    1    1    5796
0    1901    6    1    2    5804    5807
0    5808    5    1    1    5804
0    1919    6    1    2    5812    5815
0    5816    5    1    1    5812
0    5855    5    1    1    5849
0    2351    7    1    2    3751    2111
0    2366    7    3    2    3745    2105
0    2384    7    5    2    3739    2099
0    2391    7    6    2    2091    3731
0    2417    7    1    2    3725    2085
0    2431    7    2    2    3719    2335
0    2448    7    3    2    3713    2329
0    2465    7    4    2    3707    2323
0    5935    5    1    1    5929
0    2597    7    1    2    3751    2111
0    2612    7    3    2    3745    2105
0    2629    7    4    2    3739    2099
0    2635    7    5    2    3731    2091
0    2652    7    1    2    3725    2085
0    2670    7    3    2    3719    2335
0    2693    7    5    2    3713    2329
0    2715    7    6    2    3707    2323
0    6055    5    1    1    6049
0    6373    5    1    1    6367
0    6374    5    1    1    6370
0    6381    5    1    1    6375
0    6382    5    1    1    6378
0    6389    5    1    1    6383
0    6390    5    1    1    6386
0    6397    5    1    1    6391
0    6398    5    1    1    6394
0    6405    5    1    1    6399
0    6406    5    1    1    6402
0    6413    5    1    1    6407
0    6414    5    1    1    6410
0    6421    5    1    1    6415
0    6422    5    1    1    6418
0    6429    5    1    1    6423
0    6430    5    1    1    6426
0    6437    5    1    1    6431
0    6438    5    1    1    6434
0    6446    5    1    1    6442
0    3059    7    1    2    4175    3813
0    6454    5    1    1    6450
0    3068    7    1    2    4172    3810
0    6462    5    1    1    6458
0    3076    7    1    2    4169    3807
0    3079    7    1    2    4166    3804
0    6470    5    1    1    6466
0    3090    7    1    2    4163    3801
0    3099    7    1    2    4160    2175
0    3107    7    1    2    4157    2171
0    3114    7    1    2    4154    2167
0    3116    7    1    2    4151    2163
0    6502    5    1    1    6498
0    6525    5    1    1    6519
0    6526    5    1    1    6522
0    6533    5    1    1    6527
0    6534    5    1    1    6530
0    6541    5    1    1    6535
0    6542    5    1    1    6538
0    6549    5    1    1    6543
0    6550    5    1    1    6546
0    6565    5    1    1    6559
0    6566    5    1    1    6562
0    3220    5    1    1    3216
0    3292    7    1    2    4439    3838
0    3308    7    3    2    4434    3833
0    3327    7    5    2    4429    3828
0    3335    7    6    2    3821    4422
0    3362    7    1    2    4417    3816
0    3376    7    2    2    4412    2198
0    3393    7    3    2    4407    2192
0    3410    7    4    2    4402    2186
0    3425    7    5    2    4396    2179
0    6693    5    1    1    6687
0    3503    6    1    2    6687    6694
0    6701    5    1    1    6695
0    6702    5    1    1    6698
0    6709    5    1    1    6703
0    6710    5    1    1    6706
0    6728    5    1    1    6724
0    6772    5    1    1    6768
0    3853    7    1    2    4439    3838
0    3868    7    3    2    4434    3833
0    3885    7    4    2    4429    3828
0    3891    7    5    2    4422    3821
0    3908    7    1    2    4417    3816
0    3926    7    3    2    4412    2198
0    3949    7    5    2    4407    2192
0    3971    7    6    2    4402    2186
0    3979    7    7    2    4396    2179
0    7212    5    1    1    7208
0    7227    5    1    1    7221
0    7255    5    1    1    7249
0    4202    6    1    2    7249    7256
0    7263    5    1    1    7257
0    7264    5    1    1    7260
0    7272    5    1    1    7268
0    7299    5    1    1    7293
0    4225    6    1    2    7293    7300
0    7307    5    1    1    7301
0    7308    5    1    1    7304
0    7315    5    1    1    7309
0    7316    5    1    1    7312
0    4297    7    1    2    4511    2081
0    4305    7    1    2    4508    2077
0    4312    7    1    2    4505    2073
0    4314    7    1    2    4502    2069
0    4324    7    1    2    4499    2065
0    7400    5    1    1    7396
0    4333    7    1    2    4496    2316
0    7408    5    1    1    7404
0    4341    7    1    2    4493    2312
0    7416    5    1    1    7412
0    4348    7    1    2    4490    2308
0    4349    7    1    2    3686    3695
0    7431    5    1    1    7425
0    4389    7    5    2    2320    1535
0    7469    5    1    1    7463
0    4530    6    1    2    7463    7470
0    7477    5    1    1    7471
0    7478    5    1    1    7474
0    7485    5    1    1    7479
0    7486    5    1    1    7482
0    7513    5    1    1    7507
0    7514    5    1    1    7510
0    7558    5    1    1    7554
0    4932    3    2    2    917    953
0    4956    5    1    1    4952
0    4973    5    2    1    917
0    4987    5    1    1    4983
0    4997    5    1    1    4993
0    5017    5    1    1    5011
2    5099    1    877
0    5345    5    1    1    5339
0    5346    5    1    1    5342
0    5355    5    1    1    5349
0    5356    5    1    1    5352
0    5372    6    2    2    5279    5280
0    5380    6    2    2    5313    5314
0    5471    5    1    1    5465
2    5523    1    1590
0    5587    5    1    1    5581
2    5669    1    1677
2    5857    1    1841
2    5868    1    2111
2    5876    1    2105
2    5884    1    2099
2    5892    1    2091
2    5900    1    2085
2    5908    1    2335
2    5916    1    2329
2    5924    1    2323
0    5969    4    2    2    2091    3731
2    5988    1    2111
2    5996    1    2105
2    6004    1    2099
2    6012    1    2085
2    6020    1    2335
2    6028    1    2329
2    6036    1    2323
2    6044    1    2091
0    6057    4    2    2    3731    2091
2    6439    1    4175
2    6447    1    4172
2    6455    1    4169
2    6463    1    4163
2    6471    1    4160
2    6474    1    2175
2    6479    1    4157
2    6482    1    2171
2    6487    1    4154
2    6490    1    2167
2    6495    1    4166
2    6503    1    4151
2    6506    1    2163
2    6570    1    3838
2    6578    1    3833
2    6586    1    3828
2    6594    1    3821
2    6602    1    3816
2    6610    1    2198
2    6618    1    2192
2    6626    1    2186
2    6634    1    2179
0    6671    4    2    2    3821    4422
2    6721    1    2179
2    6729    1    2192
2    6732    1    2186
2    6737    1    3816
2    6740    1    2198
2    6745    1    3828
2    6748    1    3821
2    6755    1    3838
2    6758    1    3833
2    6765    1    2320
2    6773    1    2329
2    6776    1    2323
2    6781    1    2085
2    6784    1    2335
2    6789    1    2099
2    6792    1    2091
2    6799    1    2111
2    6802    1    2105
0    6832    6    2    2    6719    6720
2    6856    1    3838
2    6864    1    3833
2    6872    1    3828
2    6880    1    3816
2    6888    1    2198
2    6896    1    2192
2    6904    1    2186
2    6912    1    3821
2    6920    1    2179
0    6925    4    2    2    4422    3821
0    7041    4    2    2    4396    2179
2    7205    1    2163
2    7213    1    2171
2    7216    1    2167
2    7224    1    2175
0    7235    5    1    1    7229
0    7236    5    1    1    7232
0    7245    5    1    1    7239
0    7246    5    1    1    7242
2    7265    1    2065
2    7273    1    2073
2    7276    1    2069
2    7283    1    2081
2    7286    1    2077
0    7323    5    1    1    7317
0    7324    5    1    1    7320
0    7333    5    1    1    7327
0    7334    5    1    1    7330
2    7361    1    4511
2    7364    1    2081
2    7369    1    4508
2    7372    1    2077
2    7377    1    4505
2    7380    1    2073
2    7385    1    4499
2    7388    1    2065
2    7393    1    4496
2    7401    1    4493
2    7409    1    4490
2    7417    1    4502
2    7420    1    2069
2    7428    1    3695
0    7493    5    1    1    7487
0    7494    5    1    1    7490
0    7503    5    1    1    7497
0    7504    5    1    1    7500
2    7515    1    4493
2    7518    1    4490
2    7523    1    4499
2    7526    1    4496
2    7531    1    4505
2    7534    1    4502
2    7541    1    4511
2    7544    1    4508
2    7551    1    4151
2    7559    1    4157
2    7562    1    4154
2    7567    1    4163
2    7570    1    4160
2    7575    1    4169
2    7578    1    4166
2    7585    1    4175
2    7588    1    4172
0    1176    6    1    2    1121    1112
0    957    6    1    2    912    906
0    791    6    1    2    4881    4888
0    804    6    1    2    4889    4896
0    826    6    1    2    4897    4904
0    852    6    1    2    4905    4912
0    894    6    1    2    4921    4928
0    1025    6    1    2    5191    5198
0    1037    6    1    2    5199    5206
0    1054    6    1    2    5207    5214
0    1073    6    1    2    5215    5222
0    1092    6    1    2    5223    5230
0    1154    6    1    2    1152    1153
0    1158    6    1    2    1156    1157
0    1215    6    1    2    5250    5253
0    1224    6    1    2    5258    5261
0    1225    6    1    2    5255    5262
0    1233    6    1    2    5266    5269
0    1234    6    1    2    5263    5270
0    1238    6    1    2    5284    5287
0    1247    6    1    2    5292    5295
0    1248    6    1    2    5289    5296
0    1256    6    1    2    5300    5303
0    1257    6    1    2    5297    5304
0    1261    6    1    2    5318    5321
0    1270    6    1    2    5326    5329
0    1271    6    1    2    5323    5330
0    1279    6    1    2    5334    5337
0    1280    6    1    2    5331    5338
0    1545    6    1    2    5393    5400
0    1555    6    1    2    5401    5408
0    1572    6    1    2    5409    5416
0    1597    6    1    2    5417    5424
0    1608    6    1    2    5425    5432
0    1629    6    1    2    5433    5440
0    1654    6    1    2    5441    5448
0    1686    6    1    2    5449    5456
0    1694    6    1    2    5457    5464
0    1794    6    1    2    5745    5752
0    1804    6    1    2    5753    5760
0    1821    6    1    2    5761    5768
0    1849    6    1    2    5769    5776
0    1858    6    1    2    5777    5784
0    1868    6    1    2    5785    5792
0    1884    6    1    2    5793    5800
0    1902    6    1    2    5801    5808
0    1920    6    1    2    5809    5816
0    2954    6    1    2    6370    6373
0    2955    6    1    2    6367    6374
0    2963    6    1    2    6378    6381
0    2964    6    1    2    6375    6382
0    2971    6    1    2    6386    6389
0    2972    6    1    2    6383    6390
0    2980    6    1    2    6394    6397
0    2981    6    1    2    6391    6398
0    2990    6    1    2    6402    6405
0    2991    6    1    2    6399    6406
0    2999    6    1    2    6410    6413
0    3000    6    1    2    6407    6414
0    3007    6    1    2    6418    6421
0    3008    6    1    2    6415    6422
0    3016    6    1    2    6426    6429
0    3017    6    1    2    6423    6430
0    3019    6    1    2    6434    6437
0    3020    6    1    2    6431    6438
0    3174    6    1    2    6522    6525
0    3175    6    1    2    6519    6526
0    3184    6    1    2    6530    6533
0    3185    6    1    2    6527    6534
0    3193    6    1    2    6538    6541
0    3194    6    1    2    6535    6542
0    3201    6    1    2    6546    6549
0    3202    6    1    2    6543    6550
0    3213    6    1    2    6562    6565
0    3214    6    1    2    6559    6566
0    3227    5    1    1    3223
0    3502    6    1    2    6690    6693
0    3511    6    1    2    6698    6701
0    3512    6    1    2    6695    6702
0    3520    6    1    2    6706    6709
0    3521    6    1    2    6703    6710
0    4201    6    1    2    7252    7255
0    4210    6    1    2    7260    7263
0    4211    6    1    2    7257    7264
0    4224    6    1    2    7296    7299
0    4233    6    1    2    7304    7307
0    4234    6    1    2    7301    7308
0    4242    6    1    2    7312    7315
0    4243    6    1    2    7309    7316
0    4529    6    1    2    7466    7469
0    4538    6    1    2    7474    7477
0    4539    6    1    2    7471    7478
0    4547    6    1    2    7482    7485
0    4548    6    1    2    7479    7486
0    4552    6    1    2    7510    7513
0    4553    6    1    2    7507    7514
0    4946    5    1    1    4942
0    5347    6    1    2    5342    5345
0    5348    6    1    2    5339    5346
0    5357    6    1    2    5352    5355
0    5358    6    1    2    5349    5356
0    7237    6    1    2    7232    7235
0    7238    6    1    2    7229    7236
0    7247    6    1    2    7242    7245
0    7248    6    1    2    7239    7246
0    7325    6    1    2    7320    7323
0    7326    6    1    2    7317    7324
0    7335    6    1    2    7330    7333
0    7336    6    1    2    7327    7334
0    7495    6    1    2    7490    7493
0    7496    6    1    2    7487    7494
0    7505    6    1    2    7500    7503
0    7506    6    1    2    7497    7504
0    3244    6    1    2    3227    3220
0    792    6    7    2    790    791
0    805    6    13    2    803    804
0    827    6    15    2    825    826
0    853    6    12    2    851    852
0    895    6    6    2    893    894
0    1026    6    6    2    1024    1025
0    1038    6    9    2    1036    1037
0    1055    6    10    2    1053    1054
0    1074    6    9    2    1072    1073
0    1093    6    6    2    1091    1092
0    1155    5    1    1    1154
0    1217    6    3    2    1215    1216
0    1226    6    3    2    1224    1225
0    1235    6    2    2    1233    1234
0    1240    6    3    2    1238    1239
0    1249    6    3    2    1247    1248
0    1258    6    2    2    1256    1257
0    1263    6    3    2    1261    1262
0    1272    6    3    2    1270    1271
0    1281    6    2    2    1279    1280
0    5376    5    1    1    5372
0    5384    5    1    1    5380
0    1546    6    6    2    1544    1545
0    1556    6    10    2    1554    1555
0    1573    6    9    2    1571    1572
0    1598    6    7    2    1596    1597
0    1609    6    13    2    1607    1608
0    1630    6    15    2    1628    1629
0    1655    6    12    2    1653    1654
0    1687    6    5    2    1685    1686
0    1695    6    6    2    1693    1694
0    1795    6    6    2    1793    1794
0    1805    6    10    2    1803    1804
0    1822    6    10    2    1820    1821
0    1850    6    5    2    1848    1849
0    1859    6    6    2    1857    1858
0    1869    6    9    2    1867    1868
0    1885    6    10    2    1883    1884
0    1903    6    9    2    1901    1902
0    1921    6    6    2    1919    1920
0    5863    5    1    1    5857
0    2341    6    1    2    5868    5871
0    5872    5    1    1    5868
0    2352    6    1    2    5876    5879
0    5880    5    1    1    5876
0    2370    6    1    2    5884    5887
0    5888    5    1    1    5884
0    2398    6    1    2    5892    5895
0    5896    5    1    1    5892
0    2407    6    1    2    5900    5903
0    5904    5    1    1    5900
0    2418    6    1    2    5908    5911
0    5912    5    1    1    5908
0    2434    6    1    2    5916    5919
0    5920    5    1    1    5916
0    2452    6    1    2    5924    5927
0    5928    5    1    1    5924
0    2481    7    5    2    3682    4389
0    5975    5    1    1    5969
0    2587    6    1    2    5988    5991
0    5992    5    1    1    5988
0    2598    6    1    2    5996    5999
0    6000    5    1    1    5996
0    2616    6    1    2    6004    6007
0    6008    5    1    1    6004
0    2641    6    1    2    6012    6015
0    6016    5    1    1    6012
0    2653    6    1    2    6020    6023
0    6024    5    1    1    6020
0    2674    6    1    2    6028    6031
0    6032    5    1    1    6028
0    2699    6    1    2    6036    6039
0    6040    5    1    1    6036
0    2724    7    7    2    3682    4389
0    2732    6    1    2    6044    6047
0    6048    5    1    1    6044
0    2956    6    4    2    2954    2955
0    2965    6    3    2    2963    2964
0    2973    6    2    2    2971    2972
0    2982    6    5    2    2980    2981
0    2992    6    4    2    2990    2991
0    3001    6    3    2    2999    3000
0    3009    6    2    2    3007    3008
0    3018    6    1    2    3016    3017
0    3021    6    1    2    3019    3020
0    6445    5    1    1    6439
0    3051    6    1    2    6439    6446
0    6453    5    1    1    6447
0    3061    6    1    2    6447    6454
0    6461    5    1    1    6455
0    3070    6    1    2    6455    6462
0    6469    5    1    1    6463
0    3081    6    1    2    6463    6470
0    6477    5    1    1    6471
0    6478    5    1    1    6474
0    6485    5    1    1    6479
0    6486    5    1    1    6482
0    6493    5    1    1    6487
0    6494    5    1    1    6490
0    6501    5    1    1    6495
0    3118    6    1    2    6495    6502
0    6509    5    1    1    6503
0    6510    5    1    1    6506
0    3176    6    5    2    3174    3175
0    3186    6    4    2    3184    3185
0    3195    6    3    2    3193    3194
0    3203    6    2    2    3201    3202
0    3215    6    1    2    3213    3214
0    3281    6    1    2    6570    6573
0    6574    5    1    1    6570
0    3293    6    1    2    6578    6581
0    6582    5    1    1    6578
0    3312    6    1    2    6586    6589
0    6590    5    1    1    6586
0    3342    6    1    2    6594    6597
0    6598    5    1    1    6594
0    3351    6    1    2    6602    6605
0    6606    5    1    1    6602
0    3363    6    1    2    6610    6613
0    6614    5    1    1    6610
0    3379    6    1    2    6618    6621
0    6622    5    1    1    6618
0    3397    6    1    2    6626    6629
0    6630    5    1    1    6626
0    3415    6    1    2    6634    6637
0    6638    5    1    1    6634
0    6677    5    1    1    6671
0    3504    6    3    2    3502    3503
0    3513    6    3    2    3511    3512
0    3522    6    2    2    3520    3521
0    6727    5    1    1    6721
0    3526    6    1    2    6721    6728
0    6735    5    1    1    6729
0    6736    5    1    1    6732
0    6743    5    1    1    6737
0    6744    5    1    1    6740
0    6771    5    1    1    6765
0    3549    6    1    2    6765    6772
0    6779    5    1    1    6773
0    6780    5    1    1    6776
0    6787    5    1    1    6781
0    6788    5    1    1    6784
0    6836    5    1    1    6832
0    3843    6    1    2    6856    6859
0    6860    5    1    1    6856
0    3854    6    1    2    6864    6867
0    6868    5    1    1    6864
0    3872    6    1    2    6872    6875
0    6876    5    1    1    6872
0    3897    6    1    2    6880    6883
0    6884    5    1    1    6880
0    3909    6    1    2    6888    6891
0    6892    5    1    1    6888
0    3930    6    1    2    6896    6899
0    6900    5    1    1    6896
0    3955    6    1    2    6904    6907
0    6908    5    1    1    6904
0    3987    6    1    2    6912    6915
0    6916    5    1    1    6912
0    3995    6    1    2    6920    6923
0    6924    5    1    1    6920
0    7211    5    1    1    7205
0    4179    6    1    2    7205    7212
0    7219    5    1    1    7213
0    7220    5    1    1    7216
0    4196    6    1    2    7224    7227
0    7228    5    1    1    7224
0    4203    6    3    2    4201    4202
0    4212    6    3    2    4210    4211
0    7271    5    1    1    7265
0    4220    6    1    2    7265    7272
0    4226    6    3    2    4224    4225
0    4235    6    3    2    4233    4234
0    4244    6    2    2    4242    4243
0    7367    5    1    1    7361
0    7368    5    1    1    7364
0    7375    5    1    1    7369
0    7376    5    1    1    7372
0    7383    5    1    1    7377
0    7384    5    1    1    7380
0    7391    5    1    1    7385
0    7392    5    1    1    7388
0    7399    5    1    1    7393
0    4326    6    1    2    7393    7400
0    7407    5    1    1    7401
0    4335    6    1    2    7401    7408
0    7415    5    1    1    7409
0    4343    6    1    2    7409    7416
0    7423    5    1    1    7417
0    7424    5    1    1    7420
0    4353    6    1    2    7428    7431
0    7432    5    1    1    7428
0    4531    6    3    2    4529    4530
0    4540    6    3    2    4538    4539
0    4549    6    2    2    4547    4548
0    4554    6    3    2    4552    4553
0    7521    5    1    1    7515
0    7522    5    1    1    7518
0    7529    5    1    1    7523
0    7530    5    1    1    7526
0    7557    5    1    1    7551
0    4576    6    1    2    7551    7558
0    7565    5    1    1    7559
0    7566    5    1    1    7562
0    7573    5    1    1    7567
0    7574    5    1    1    7570
0    4936    5    1    1    4932
0    4937    6    1    2    4932    4935
0    4977    5    1    1    4973
0    4978    6    1    2    4973    4976
0    5105    5    1    1    5099
0    5359    6    2    2    5357    5358
0    5362    6    2    2    5347    5348
0    5529    5    1    1    5523
0    5675    5    1    1    5669
2    5932    1    4389
2    5977    1    2391
2    6052    1    4389
0    6063    5    1    1    6057
2    6115    1    2635
0    6173    4    2    2    3682    4389
2    6679    1    3335
0    6751    5    1    1    6745
0    6752    5    1    1    6748
0    6761    5    1    1    6755
0    6762    5    1    1    6758
0    6795    5    1    1    6789
0    6796    5    1    1    6792
0    6805    5    1    1    6799
0    6806    5    1    1    6802
0    6931    5    1    1    6925
2    6983    1    3891
0    7047    5    1    1    7041
2    7129    1    3979
0    7279    5    1    1    7273
0    7280    5    1    1    7276
0    7289    5    1    1    7283
0    7290    5    1    1    7286
0    7337    6    2    2    7247    7248
0    7340    6    2    2    7237    7238
0    7353    6    2    2    7335    7336
0    7356    6    2    2    7325    7326
0    7537    5    1    1    7531
0    7538    5    1    1    7534
0    7547    5    1    1    7541
0    7548    5    1    1    7544
0    7581    5    1    1    7575
0    7582    5    1    1    7578
0    7591    5    1    1    7585
0    7592    5    1    1    7588
0    7595    6    2    2    7505    7506
0    7598    6    2    2    7495    7496
0    2342    6    1    2    5865    5872
0    2353    6    1    2    5873    5880
0    2371    6    1    2    5881    5888
0    2399    6    1    2    5889    5896
0    2408    6    1    2    5897    5904
0    2419    6    1    2    5905    5912
0    2435    6    1    2    5913    5920
0    2453    6    1    2    5921    5928
0    2588    6    1    2    5985    5992
0    2599    6    1    2    5993    6000
0    2617    6    1    2    6001    6008
0    2642    6    1    2    6009    6016
0    2654    6    1    2    6017    6024
0    2675    6    1    2    6025    6032
0    2700    6    1    2    6033    6040
0    2733    6    1    2    6041    6048
0    3050    6    1    2    6442    6445
0    3060    6    1    2    6450    6453
0    3069    6    1    2    6458    6461
0    3080    6    1    2    6466    6469
0    3091    6    1    2    6474    6477
0    3092    6    1    2    6471    6478
0    3100    6    1    2    6482    6485
0    3101    6    1    2    6479    6486
0    3108    6    1    2    6490    6493
0    3109    6    1    2    6487    6494
0    3117    6    1    2    6498    6501
0    3120    6    1    2    6506    6509
0    3121    6    1    2    6503    6510
0    3282    6    1    2    6567    6574
0    3294    6    1    2    6575    6582
0    3313    6    1    2    6583    6590
0    3343    6    1    2    6591    6598
0    3352    6    1    2    6599    6606
0    3364    6    1    2    6607    6614
0    3380    6    1    2    6615    6622
0    3398    6    1    2    6623    6630
0    3416    6    1    2    6631    6638
0    3525    6    1    2    6724    6727
0    3534    6    1    2    6732    6735
0    3535    6    1    2    6729    6736
0    3543    6    1    2    6740    6743
0    3544    6    1    2    6737    6744
0    3548    6    1    2    6768    6771
0    3557    6    1    2    6776    6779
0    3558    6    1    2    6773    6780
0    3566    6    1    2    6784    6787
0    3567    6    1    2    6781    6788
0    3844    6    1    2    6853    6860
0    3855    6    1    2    6861    6868
0    3873    6    1    2    6869    6876
0    3898    6    1    2    6877    6884
0    3910    6    1    2    6885    6892
0    3931    6    1    2    6893    6900
0    3956    6    1    2    6901    6908
0    3988    6    1    2    6909    6916
0    3996    6    1    2    6917    6924
0    4178    6    1    2    7208    7211
0    4187    6    1    2    7216    7219
0    4188    6    1    2    7213    7220
0    4197    6    1    2    7221    7228
0    4219    6    1    2    7268    7271
0    4289    6    1    2    7364    7367
0    4290    6    1    2    7361    7368
0    4298    6    1    2    7372    7375
0    4299    6    1    2    7369    7376
0    4306    6    1    2    7380    7383
0    4307    6    1    2    7377    7384
0    4315    6    1    2    7388    7391
0    4316    6    1    2    7385    7392
0    4325    6    1    2    7396    7399
0    4334    6    1    2    7404    7407
0    4342    6    1    2    7412    7415
0    4350    6    1    2    7420    7423
0    4351    6    1    2    7417    7424
0    4354    6    1    2    7425    7432
0    4561    6    1    2    7518    7521
0    4562    6    1    2    7515    7522
0    4570    6    1    2    7526    7529
0    4571    6    1    2    7523    7530
0    4575    6    1    2    7554    7557
0    4584    6    1    2    7562    7565
0    4585    6    1    2    7559    7566
0    4593    6    1    2    7570    7573
0    4594    6    1    2    7567    7574
0    4938    6    1    2    4929    4936
0    4979    6    1    2    4970    4977
0    6753    6    1    2    6748    6751
0    6754    6    1    2    6745    6752
0    6763    6    1    2    6758    6761
0    6764    6    1    2    6755    6762
0    6797    6    1    2    6792    6795
0    6798    6    1    2    6789    6796
0    6807    6    1    2    6802    6805
0    6808    6    1    2    6799    6806
0    7281    6    1    2    7276    7279
0    7282    6    1    2    7273    7280
0    7291    6    1    2    7286    7289
0    7292    6    1    2    7283    7290
0    7539    6    1    2    7534    7537
0    7540    6    1    2    7531    7538
0    7549    6    1    2    7544    7547
0    7550    6    1    2    7541    7548
0    7583    6    1    2    7578    7581
0    7584    6    1    2    7575    7582
0    7593    6    1    2    7588    7591
0    7594    6    1    2    7585    7592
0    1856    5    1    1    1850
0    920    7    3    5    895    853    827    805    792
0    925    7    1    2    792    821
0    926    7    1    3    805    792    845
0    927    7    1    4    827    792    868    805
0    928    7    1    5    853    827    792    877    805
0    937    7    1    2    805    845
0    938    7    1    3    827    868    805
0    939    7    1    4    853    827    877    805
0    940    7    1    4    895    827    805    853
0    941    7    1    2    805    845
0    942    7    1    3    827    868    805
0    943    7    1    4    853    827    877    805
0    944    7    1    2    827    868
0    945    7    1    3    853    827    877
0    946    7    1    3    895    827    853
0    947    7    1    2    827    868
0    948    7    1    3    853    827    877
0    949    7    1    2    853    877
0    956    7    1    2    895    853
0    1122    7    2    5    1038    1093    1055    1026    1074
0    1125    7    1    2    1026    1050
0    1126    7    1    3    1038    1026    1068
0    1127    7    1    4    1055    1026    1086    1038
0    1128    7    1    5    1074    1055    1026    1102    1038
0    1132    7    1    2    1038    1068
0    1133    7    1    3    1055    1086    1038
0    1134    7    1    4    1074    1055    1102    1038
0    1137    7    1    2    1086    1055
0    1138    7    1    3    1074    1055    1102
0    1141    7    1    2    1074    1102
0    1221    5    2    1    1217
0    1230    5    2    1    1226
0    1244    5    2    1    1240
0    1253    5    2    1    1249
0    1267    5    2    1    1263
0    1276    5    2    1    1272
2    1284    1    1235
2    1288    1    1235
2    1292    1    1258
2    1296    1    1258
2    1300    1    1281
2    1304    1    1281
0    1702    7    2    4    1687    1573    1556    1546
0    1705    7    1    2    1546    1567
0    1706    7    1    3    1556    1546    1584
0    1707    7    1    4    1573    1546    1590    1556
0    1709    7    1    2    1556    1584
0    1710    7    1    3    1573    1590    1556
0    1711    7    1    3    1687    1573    1556
0    1712    7    1    2    1556    1584
0    1713    7    1    3    1573    1590    1556
0    1714    7    1    2    1573    1590
0    1718    7    2    5    1695    1655    1630    1609    1598
0    1722    7    1    2    1598    1624
0    1723    7    1    3    1609    1598    1647
0    1724    7    1    4    1630    1598    1669    1609
0    1725    7    1    5    1655    1630    1598    1677    1609
0    1733    7    1    2    1609    1647
0    1734    7    1    3    1630    1669    1609
0    1735    7    1    4    1655    1630    1677    1609
0    1736    7    1    4    1695    1630    1609    1655
0    1737    7    1    2    1609    1647
0    1738    7    1    3    1630    1669    1609
0    1739    7    1    4    1655    1630    1677    1609
0    1740    7    1    2    1630    1669
0    1741    7    1    3    1655    1630    1677
0    1742    7    1    3    1695    1630    1655
0    1743    7    1    2    1630    1669
0    1744    7    1    3    1655    1630    1677
0    1745    7    1    2    1655    1677
0    1749    7    1    2    1687    1573
0    1750    7    1    2    1695    1655
0    1935    7    2    4    1805    1850    1822    1795
0    1938    7    1    2    1795    1816
0    1939    7    1    3    1805    1795    1834
0    1940    7    1    4    1822    1795    1841    1805
0    1942    7    1    2    1805    1834
0    1943    7    1    3    1822    1841    1805
0    1944    7    1    3    1850    1822    1805
0    1945    7    1    2    1805    1834
0    1946    7    1    3    1841    1822    1805
0    1947    7    1    2    1822    1841
0    1948    7    1    2    1850    1822
0    1949    7    1    2    1822    1841
0    1950    7    2    5    1869    1921    1885    1859    1903
0    1953    7    1    2    1859    1880
0    1954    7    1    3    1869    1859    1897
0    1955    7    1    4    1885    1859    1914    1869
0    1956    7    1    5    1903    1885    1859    1929    1869
0    1960    7    1    2    1869    1897
0    1961    7    1    3    1885    1914    1869
0    1962    7    1    4    1903    1885    1929    1869
0    1965    7    1    2    1914    1885
0    1966    7    1    3    1903    1885    1929
0    1969    7    1    2    1903    1929
0    2343    6    6    2    2341    2342
0    2354    6    10    2    2352    2353
0    2372    6    10    2    2370    2371
0    2400    6    5    2    2398    2399
0    2409    6    6    2    2407    2408
0    2420    6    9    2    2418    2419
0    2436    6    10    2    2434    2435
0    2454    6    9    2    2452    2453
0    2470    6    1    2    5932    5935
0    5936    5    1    1    5932
0    5983    5    1    1    5977
0    2589    6    6    2    2587    2588
0    2600    6    10    2    2598    2599
0    2618    6    9    2    2616    2617
0    2643    6    7    2    2641    2642
0    2655    6    13    2    2653    2654
0    2676    6    15    2    2674    2675
0    2701    6    12    2    2699    2700
0    2734    6    5    2    2732    2733
0    2740    6    1    2    6052    6055
0    6056    5    1    1    6052
0    3022    7    2    4    3018    2973    2965    2956
0    3025    7    1    2    2956    2970
0    3026    7    1    3    2965    2956    2977
0    3027    7    1    4    2973    2956    2979    2965
0    3029    7    1    5    3021    3009    3001    2992    2982
0    3030    7    1    2    2982    2998
0    3031    7    1    3    2992    2982    3006
0    3032    7    1    4    3001    2982    3013    2992
0    3033    7    1    5    3009    3001    2982    3015    2992
0    3052    6    4    2    3050    3051
0    3062    6    3    2    3060    3061
0    3071    6    2    2    3069    3070
0    3082    6    5    2    3080    3081
0    3093    6    4    2    3091    3092
0    3102    6    3    2    3100    3101
0    3110    6    2    2    3108    3109
0    3119    6    1    2    3117    3118
0    3122    6    1    2    3120    3121
0    3228    7    2    5    3215    3203    3195    3186    3176
0    3231    7    1    2    3176    3192
0    3232    7    1    3    3186    3176    3200
0    3233    7    1    4    3195    3176    3207    3186
0    3234    7    1    5    3203    3195    3176    3209    3186
0    3283    6    6    2    3281    3282
0    3295    6    10    2    3293    3294
0    3314    6    10    2    3312    3313
0    3344    6    5    2    3342    3343
0    3353    6    6    2    3351    3352
0    3365    6    9    2    3363    3364
0    3381    6    10    2    3379    3380
0    3399    6    9    2    3397    3398
0    3417    6    6    2    3415    3416
0    6685    5    1    1    6679
0    3508    5    2    1    3504
0    3517    5    2    1    3513
0    3527    6    3    2    3525    3526
0    3536    6    3    2    3534    3535
0    3545    6    2    2    3543    3544
0    3550    6    3    2    3548    3549
0    3559    6    3    2    3557    3558
0    3568    6    2    2    3566    3567
2    3571    1    3522
2    3575    1    3522
0    3845    6    6    2    3843    3844
0    3856    6    10    2    3854    3855
0    3874    6    9    2    3872    3873
0    3899    6    7    2    3897    3898
0    3911    6    13    2    3909    3910
0    3932    6    15    2    3930    3931
0    3957    6    12    2    3955    3956
0    3989    6    5    2    3987    3988
0    3997    6    6    2    3995    3996
0    4180    6    3    2    4178    4179
0    4189    6    3    2    4187    4188
0    4198    6    2    2    4196    4197
0    4207    5    2    1    4203
0    4216    5    2    1    4212
0    4221    6    2    2    4219    4220
0    4230    5    2    1    4226
0    4239    5    2    1    4235
2    4263    1    4244
2    4267    1    4244
0    4291    6    4    2    4289    4290
0    4300    6    3    2    4298    4299
0    4308    6    2    2    4306    4307
0    4317    6    5    2    4315    4316
0    4327    6    4    2    4325    4326
0    4336    6    3    2    4334    4335
0    4344    6    2    2    4342    4343
0    4352    6    1    2    4350    4351
0    4355    6    1    2    4353    4354
0    4535    5    2    1    4531
0    4544    5    2    1    4540
0    4558    5    2    1    4554
0    4563    6    3    2    4561    4562
0    4572    6    2    2    4570    4571
0    4577    6    3    2    4575    4576
0    4586    6    3    2    4584    4585
0    4595    6    2    2    4593    4594
2    4598    1    4549
2    4602    1    4549
2    4716    1    1921
2    4724    1    1859
2    4732    1    1869
2    4740    1    1885
2    4748    1    1903
2    4756    1    1093
2    4764    1    1026
2    4772    1    1038
2    4780    1    1055
2    4788    1    1074
0    4939    6    2    2    4937    4938
0    4980    6    2    2    4978    4979
2    5044    1    895
2    5054    1    853
2    5064    1    792
2    5074    1    827
2    5084    1    805
2    5094    1    805
2    5132    1    895
2    5142    1    853
2    5152    1    792
2    5162    1    827
0    5365    5    1    1    5359
0    5366    5    1    1    5362
2    5488    1    1687
2    5498    1    1573
2    5508    1    1546
2    5518    1    1556
2    5546    1    1687
2    5556    1    1573
2    5566    1    1546
2    5576    1    1556
2    5614    1    1695
2    5624    1    1655
2    5634    1    1598
2    5644    1    1630
2    5654    1    1609
2    5664    1    1609
2    5702    1    1695
2    5712    1    1655
2    5722    1    1598
2    5732    1    1630
2    5820    1    1795
2    5828    1    1795
2    5836    1    1805
2    5844    1    1805
2    5852    1    1822
2    5860    1    1822
0    6121    5    1    1    6115
0    6179    5    1    1    6173
2    6261    1    2724
0    7359    5    1    1    7353
0    7360    5    1    1    7356
0    7343    5    1    1    7337
0    7344    5    1    1    7340
0    6809    6    2    2    6763    6764
0    6812    6    2    2    6753    6754
0    6819    6    2    2    6807    6808
0    6822    6    2    2    6797    6798
0    6989    5    1    1    6983
0    7135    5    1    1    7129
0    7345    6    2    2    7291    7292
0    7348    6    2    2    7281    7282
0    7601    5    1    1    7595
0    7602    5    1    1    7598
0    7603    6    2    2    7549    7550
0    7606    6    2    2    7539    7540
0    7611    6    2    2    7593    7594
0    7614    6    2    2    7583    7584
0    929    3    3    5    802    925    926    927    928
0    950    3    2    2    868    949
0    1129    3    2    5    1035    1125    1126    1127    1128
0    1708    3    1    4    1553    1705    1706    1707
0    1715    3    2    2    1584    1714
0    1726    3    3    5    1606    1722    1723    1724    1725
0    1746    3    2    2    1669    1745
0    1941    3    1    4    1802    1938    1939    1940
0    1957    3    2    5    1866    1953    1954    1955    1956
0    2471    6    1    2    5929    5936
0    2741    6    1    2    6049    6056
0    3028    3    1    4    2962    3025    3026    3027
0    3034    3    1    5    2989    3030    3031    3032    3033
0    3235    3    2    5    3183    3231    3232    3233    3234
0    5014    3    2    4    845    944    945    946
0    5034    3    2    5    821    937    938    939    940
0    5102    4    2    3    845    947    948
0    5122    4    2    4    821    941    942    943
0    5367    6    1    2    5362    5365
0    5368    6    1    2    5359    5366
0    5478    3    2    4    1567    1709    1710    1711
0    5536    4    2    3    1567    1712    1713
0    5584    3    2    4    1647    1740    1741    1742
0    5604    3    2    5    1624    1733    1734    1735    1736
0    5672    4    2    3    1647    1743    1744
0    5692    4    2    4    1624    1737    1738    1739
0    5817    3    2    4    1816    1942    1943    1944
0    5825    4    2    3    1816    1945    1946
0    5833    3    2    3    1834    1947    1948
0    5841    4    2    2    1834    1949
0    6340    6    1    2    7356    7359
0    6341    6    1    2    7353    7360
0    6350    6    1    2    7340    7343
0    6351    6    1    2    7337    7344
0    7436    6    1    2    7598    7601
0    7437    6    1    2    7595    7602
0    4720    5    1    1    4716
0    4728    5    1    1    4724
0    4736    5    1    1    4732
0    4744    5    1    1    4740
0    4752    5    1    1    4748
0    4760    5    1    1    4756
0    4768    5    1    1    4764
0    4776    5    1    1    4772
0    4784    5    1    1    4780
0    4792    5    1    1    4788
0    3350    5    1    1    3344
0    2406    5    1    1    2400
0    924    5    1    1    920
0    5088    5    1    1    5084
0    5098    5    1    1    5094
0    997    7    4    2    902    920
0    1146    7    4    2    1108    1122
0    1287    5    1    1    1284
0    1291    5    1    1    1288
0    1295    5    1    1    1292
0    1299    5    1    1    1296
0    1303    5    1    1    1300
0    1307    5    1    1    1304
0    1309    7    1    3    1226    1217    1284
0    1312    7    1    3    1230    1221    1288
0    1315    7    1    3    1249    1240    1292
0    1318    7    1    3    1253    1244    1296
0    1321    7    1    3    1272    1263    1300
0    1324    7    1    3    1276    1267    1304
0    1721    5    1    1    1718
0    5522    5    1    1    5518
0    5580    5    1    1    5576
0    5658    5    1    1    5654
0    5668    5    1    1    5664
0    1788    7    6    2    1702    1718
0    1974    7    6    2    1935    1950
0    5824    5    1    1    5820
0    5832    5    1    1    5828
0    5840    5    1    1    5836
0    5848    5    1    1    5844
0    1999    6    1    2    5852    5855
0    5856    5    1    1    5852
0    2003    6    1    2    5860    5863
0    5864    5    1    1    5860
0    2472    6    6    2    2470    2471
0    2487    7    3    4    2354    2400    2372    2343
0    2492    7    1    2    2343    2366
0    2493    7    1    3    2354    2343    2384
0    2494    7    1    4    2372    2343    2391    2354
0    2500    7    1    2    2354    2384
0    2501    7    1    3    2372    2391    2354
0    2502    7    1    3    2400    2372    2354
0    2503    7    1    2    2354    2384
0    2504    7    1    3    2391    2372    2354
0    2505    7    1    2    2372    2391
0    2506    7    1    2    2400    2372
0    2507    7    1    2    2372    2391
0    2511    7    1    2    2409    2431
0    2512    7    1    3    2420    2409    2448
0    2513    7    1    4    2436    2409    2465    2420
0    2514    7    1    5    2454    2436    2409    2481    2420
0    2518    7    1    2    2420    2448
0    2519    7    1    3    2436    2465    2420
0    2520    7    1    4    2454    2436    2481    2420
0    2523    7    1    2    2465    2436
0    2524    7    1    3    2454    2436    2481
0    2527    7    1    2    2454    2481
0    2742    6    6    2    2740    2741
0    2749    7    3    4    2734    2618    2600    2589
0    2754    7    1    2    2589    2612
0    2755    7    1    3    2600    2589    2629
0    2756    7    1    4    2618    2589    2635    2600
0    2762    7    1    2    2600    2629
0    2763    7    1    3    2618    2635    2600
0    2764    7    1    3    2734    2618    2600
0    2765    7    1    2    2600    2629
0    2766    7    1    3    2618    2635    2600
0    2767    7    1    2    2618    2635
0    2776    7    1    2    2643    2670
0    2777    7    1    3    2655    2643    2693
0    2778    7    1    4    2676    2643    2715    2655
0    2779    7    1    5    2701    2676    2643    2724    2655
0    2788    7    1    2    2655    2693
0    2789    7    1    3    2676    2715    2655
0    2790    7    1    4    2701    2676    2724    2655
0    2792    7    1    2    2655    2693
0    2793    7    1    3    2676    2715    2655
0    2794    7    1    4    2701    2676    2724    2655
0    2795    7    1    2    2676    2715
0    2796    7    1    3    2701    2676    2724
0    2798    7    1    2    2676    2715
0    2799    7    1    3    2701    2676    2724
0    2800    7    1    2    2701    2724
0    2804    7    1    2    2734    2618
0    3035    7    9    2    3022    3029
0    3045    7    1    2    3022    3034
0    3123    7    3    4    3119    3071    3062    3052
0    3128    7    1    2    3052    3068
0    3129    7    1    3    3062    3052    3076
0    3130    7    1    4    3071    3052    3079    3062
0    3136    7    2    5    3122    3110    3102    3093    3082
0    3139    7    1    2    3082    3099
0    3140    7    1    3    3093    3082    3107
0    3141    7    1    4    3102    3082    3114    3093
0    3142    7    1    5    3110    3102    3082    3116    3093
0    3249    7    8    2    3216    3228
0    3431    7    2    4    3295    3344    3314    3283
0    3434    7    1    2    3283    3308
0    3435    7    1    3    3295    3283    3327
0    3436    7    1    4    3314    3283    3335    3295
0    3438    7    1    2    3295    3327
0    3439    7    1    3    3314    3335    3295
0    3440    7    1    3    3344    3314    3295
0    3441    7    1    2    3295    3327
0    3442    7    1    3    3335    3314    3295
0    3443    7    1    2    3314    3335
0    3444    7    1    2    3344    3314
0    3445    7    1    2    3314    3335
0    3446    7    2    5    3365    3417    3381    3353    3399
0    3449    7    1    2    3353    3376
0    3450    7    1    3    3365    3353    3393
0    3451    7    1    4    3381    3353    3410    3365
0    3452    7    1    5    3399    3381    3353    3425    3365
0    3456    7    1    2    3365    3393
0    3457    7    1    3    3381    3410    3365
0    3458    7    1    4    3399    3381    3425    3365
0    3460    7    1    2    3410    3381
0    3461    7    1    3    3399    3381    3425
0    3463    7    1    2    3399    3425
0    3531    5    2    1    3527
0    3540    5    2    1    3536
0    3554    5    2    1    3550
0    3563    5    2    1    3559
0    3574    5    1    1    3571
0    3578    5    1    1    3575
2    3579    1    3545
2    3583    1    3545
2    3587    1    3568
2    3591    1    3568
0    3596    7    1    3    3513    3504    3571
0    3599    7    1    3    3517    3508    3575
0    4004    7    2    4    3989    3874    3856    3845
0    4007    7    1    2    3845    3868
0    4008    7    1    3    3856    3845    3885
0    4009    7    1    4    3874    3845    3891    3856
0    4011    7    1    2    3856    3885
0    4012    7    1    3    3874    3891    3856
0    4013    7    1    3    3989    3874    3856
0    4014    7    1    2    3856    3885
0    4015    7    1    3    3874    3891    3856
0    4016    7    1    2    3874    3891
0    4020    7    2    5    3997    3957    3932    3911    3899
0    4024    7    1    2    3899    3926
0    4025    7    1    3    3911    3899    3949
0    4026    7    1    4    3932    3899    3971    3911
0    4027    7    1    5    3957    3932    3899    3979    3911
0    4035    7    1    2    3911    3949
0    4036    7    1    3    3932    3971    3911
0    4037    7    1    4    3957    3932    3979    3911
0    4038    7    1    4    3997    3932    3911    3957
0    4039    7    1    2    3911    3949
0    4040    7    1    3    3932    3971    3911
0    4041    7    1    4    3957    3932    3979    3911
0    4042    7    1    2    3932    3971
0    4043    7    1    3    3957    3932    3979
0    4044    7    1    3    3997    3932    3957
0    4045    7    1    2    3932    3971
0    4046    7    1    3    3957    3932    3979
0    4047    7    1    2    3957    3979
0    4051    7    1    2    3989    3874
0    4052    7    1    2    3997    3957
0    4184    5    2    1    4180
0    4193    5    2    1    4189
2    4247    1    4198
2    4251    1    4198
2    4255    1    4221
2    4259    1    4221
0    4266    5    1    1    4263
0    4270    5    1    1    4267
0    4284    7    1    3    4235    4226    4263
0    4287    7    1    3    4239    4230    4267
0    4356    7    3    4    4352    4308    4300    4291
0    4361    7    1    2    4291    4305
0    4362    7    1    3    4300    4291    4312
0    4363    7    1    4    4308    4291    4314    4300
0    4369    7    2    5    4355    4344    4336    4327    4317
0    4372    7    1    2    4317    4333
0    4373    7    1    3    4327    4317    4341
0    4374    7    1    4    4336    4317    4348    4327
0    4375    7    1    5    4344    4336    4317    4349    4327
0    4567    5    2    1    4563
0    4581    5    2    1    4577
0    4590    5    2    1    4586
0    4601    5    1    1    4598
0    4605    5    1    1    4602
2    4606    1    4572
2    4610    1    4572
2    4614    1    4595
2    4618    1    4595
0    4623    7    1    3    4540    4531    4598
0    4626    7    1    3    4544    4535    4602
2    4796    1    3417
2    4804    1    3353
2    4812    1    3365
2    4820    1    3381
2    4828    1    3399
2    4844    1    2409
2    4852    1    2420
2    4860    1    2436
2    4868    1    2454
0    4945    5    1    1    4939
0    4948    6    1    2    4939    4946
0    4986    5    1    1    4980
0    4989    6    1    2    4980    4987
0    5048    5    1    1    5044
0    5058    5    1    1    5054
0    5068    5    1    1    5064
0    5078    5    1    1    5074
0    5166    5    1    1    5162
0    5136    5    1    1    5132
0    5146    5    1    1    5142
0    5156    5    1    1    5152
0    5388    6    2    2    5367    5368
0    5492    5    1    1    5488
0    5502    5    1    1    5498
0    5512    5    1    1    5508
0    5550    5    1    1    5546
0    5560    5    1    1    5556
0    5570    5    1    1    5566
0    5618    5    1    1    5614
0    5628    5    1    1    5624
0    5638    5    1    1    5634
0    5648    5    1    1    5644
0    5736    5    1    1    5732
0    5706    5    1    1    5702
0    5716    5    1    1    5712
0    5726    5    1    1    5722
2    5940    1    2343
2    5948    1    2343
2    5956    1    2354
2    5964    1    2354
2    5972    1    2372
2    5980    1    2372
2    6080    1    2734
2    6090    1    2618
2    6100    1    2589
2    6110    1    2600
2    6138    1    2734
2    6148    1    2618
2    6158    1    2589
2    6168    1    2600
2    6216    1    2701
2    6226    1    2643
2    6236    1    2676
2    6246    1    2655
2    6256    1    2655
0    6267    5    1    1    6261
2    6304    1    2701
2    6314    1    2643
2    6324    1    2676
0    6342    6    2    2    6340    6341
0    6352    6    2    2    6350    6351
0    7351    5    1    1    7345
0    7352    5    1    1    7348
2    6642    1    3283
2    6650    1    3283
2    6658    1    3295
2    6666    1    3295
2    6674    1    3314
2    6682    1    3314
0    6815    5    1    1    6809
0    6816    5    1    1    6812
0    6825    5    1    1    6819
0    6826    5    1    1    6822
2    6948    1    3989
2    6958    1    3874
2    6968    1    3845
2    6978    1    3856
2    7006    1    3989
2    7016    1    3874
2    7026    1    3845
2    7036    1    3856
2    7074    1    3997
2    7084    1    3957
2    7094    1    3899
2    7104    1    3932
2    7114    1    3911
2    7124    1    3911
2    7162    1    3997
2    7172    1    3957
2    7182    1    3899
2    7192    1    3932
0    7438    6    2    2    7436    7437
0    7617    5    1    1    7611
0    7618    5    1    1    7614
0    7609    5    1    1    7603
0    7610    5    1    1    7606
0    1151    7    1    2    1129    1108
0    1002    7    1    2    902    929
0    933    5    3    1    929
0    1308    7    1    3    1221    1226    1287
0    1311    7    1    3    1217    1230    1291
0    1314    7    1    3    1244    1249    1295
0    1317    7    1    3    1240    1253    1299
0    1320    7    1    3    1267    1272    1303
0    1323    7    1    3    1263    1276    1307
0    1730    5    2    1    1726
0    1789    7    1    2    1702    1726
0    1981    7    1    2    1957    1935
0    5823    5    1    1    5817
0    1986    6    1    2    5817    5824
0    5831    5    1    1    5825
0    1989    6    1    2    5825    5832
0    5839    5    1    1    5833
0    1993    6    1    2    5833    5840
0    5847    5    1    1    5841
0    1996    6    1    2    5841    5848
0    2000    6    1    2    5849    5856
0    2004    6    1    2    5857    5864
0    2495    3    3    4    2351    2492    2493    2494
0    2515    3    2    5    2417    2511    2512    2513    2514
0    2757    3    3    4    2597    2754    2755    2756
0    2768    3    2    2    2629    2767
0    2780    3    3    5    2652    2776    2777    2778    2779
0    2801    3    2    2    2715    2800
0    3046    3    3    2    3028    3045
0    3131    3    3    4    3059    3128    3129    3130
0    3143    3    2    5    3090    3139    3140    3141    3142
0    3238    5    1    1    3235
0    3258    7    1    2    3216    3235
0    3437    3    1    4    3292    3434    3435    3436
0    3453    3    2    5    3362    3449    3450    3451    3452
0    3595    7    1    3    3508    3513    3574
0    3598    7    1    3    3504    3517    3578
0    4010    3    1    4    3853    4007    4008    4009
0    4017    3    2    2    3885    4016
0    4028    3    3    5    3908    4024    4025    4026    4027
0    4048    3    2    2    3971    4047
0    4283    7    1    3    4230    4235    4266
0    4286    7    1    3    4226    4239    4270
0    4364    3    3    4    4297    4361    4362    4363
0    4376    3    2    5    4324    4372    4373    4374    4375
0    4622    7    1    3    4535    4540    4601
0    4625    7    1    3    4531    4544    4605
0    4947    6    1    2    4942    4945
0    4988    6    1    2    4983    4986
0    5018    5    1    1    5014
0    5019    6    1    2    5014    5017
0    5024    3    2    2    950    956
0    5038    5    1    1    5034
0    5106    5    1    1    5102
0    5107    6    1    2    5102    5105
0    5112    5    2    1    950
0    5126    5    1    1    5122
0    5468    3    2    2    1715    1749
0    5482    5    1    1    5478
0    5526    5    2    1    1715
0    5540    5    1    1    5536
0    5588    5    1    1    5584
0    5589    6    1    2    5584    5587
0    5594    3    2    2    1746    1750
0    5608    5    1    1    5604
0    5676    5    1    1    5672
0    5677    6    1    2    5672    5675
0    5682    5    2    1    1746
0    5696    5    1    1    5692
0    5937    3    2    4    2366    2500    2501    2502
0    5945    4    2    3    2366    2503    2504
0    5953    3    2    3    2384    2505    2506
0    5961    4    2    2    2384    2507
0    6070    3    2    4    2612    2762    2763    2764
0    6128    4    2    3    2612    2765    2766
0    6264    4    2    3    2693    2798    2799
0    6284    4    2    4    2670    2792    2793    2794
0    6360    6    1    2    7348    7351
0    6361    6    1    2    7345    7352
0    6639    3    2    4    3308    3438    3439    3440
0    6647    4    2    3    3308    3441    3442
0    6655    3    2    3    3327    3443    3444
0    6663    4    2    2    3327    3445
0    6817    6    1    2    6812    6815
0    6818    6    1    2    6809    6816
0    6827    6    1    2    6822    6825
0    6828    6    1    2    6819    6826
0    6938    3    2    4    3868    4011    4012    4013
0    6996    4    2    3    3868    4014    4015
0    7044    3    2    4    3949    4042    4043    4044
0    7064    3    2    5    3926    4035    4036    4037    4038
0    7132    4    2    3    3949    4045    4046
0    7152    4    2    4    3926    4039    4040    4041
0    7446    6    1    2    7614    7617
0    7447    6    1    2    7611    7618
0    7456    6    1    2    7606    7609
0    7457    6    1    2    7603    7610
0    241    3    1    2    1117    1151
0    265    3    1    2    908    1002
0    2005    6    1    2    2003    2004
0    4800    5    1    1    4796
0    4808    5    1    1    4804
0    4816    5    1    1    4812
0    4824    5    1    1    4820
0    4832    5    1    1    4828
0    4848    5    1    1    4844
0    4856    5    1    1    4852
0    4864    5    1    1    4860
0    4872    5    1    1    4868
0    1310    4    1    2    1308    1309
0    1313    4    1    2    1311    1312
0    1316    4    1    2    1314    1315
0    1319    4    1    2    1317    1318
0    1322    4    1    2    1320    1321
0    1325    4    1    2    1323    1324
0    5392    5    1    1    5388
0    1790    3    2    2    1708    1789
0    1982    3    2    2    1941    1981
0    1985    6    1    2    5820    5823
0    1988    6    1    2    5828    5831
0    1992    6    1    2    5836    5839
0    1995    6    1    2    5844    5847
0    2001    6    1    2    1999    2000
0    2491    5    1    1    2487
0    2508    7    2    5    2420    2472    2436    2409    2454
0    2522    7    1    5    4526    2472    2436    2454    2420
0    2526    7    1    4    4526    2472    2436    2454
0    2529    7    1    3    4526    2472    2454
0    2531    7    1    2    4526    2472
0    5944    5    1    1    5940
0    5952    5    1    1    5948
0    5960    5    1    1    5956
0    5968    5    1    1    5964
0    2555    6    1    2    5972    5975
0    5976    5    1    1    5972
0    2559    6    1    2    5980    5983
0    5984    5    1    1    5980
0    2753    5    1    1    2749
0    2771    7    3    5    2742    2701    2676    2655    2643
0    2791    7    1    4    2742    2676    2655    2701
0    2797    7    1    3    2742    2676    2701
0    2807    7    1    2    2742    2701
0    6114    5    1    1    6110
0    6172    5    1    1    6168
0    6250    5    1    1    6246
0    6260    5    1    1    6256
0    6346    5    1    1    6342
0    6356    5    1    1    6352
0    3127    5    1    1    3123
0    3156    7    6    2    3123    3136
0    3259    3    2    2    3223    3258
0    3466    7    6    2    3431    3446
0    6646    5    1    1    6642
0    6654    5    1    1    6650
0    6662    5    1    1    6658
0    6670    5    1    1    6666
0    3483    6    1    2    6674    6677
0    6678    5    1    1    6674
0    3487    6    1    2    6682    6685
0    6686    5    1    1    6682
0    3582    5    1    1    3579
0    3586    5    1    1    3583
0    3590    5    1    1    3587
0    3594    5    1    1    3591
0    3597    4    1    2    3595    3596
0    3600    4    1    2    3598    3599
0    3602    7    1    3    3536    3527    3579
0    3605    7    1    3    3540    3531    3583
0    3608    7    1    3    3559    3550    3587
0    3611    7    1    3    3563    3554    3591
0    4023    5    1    1    4020
0    6982    5    1    1    6978
0    7040    5    1    1    7036
0    7118    5    1    1    7114
0    7128    5    1    1    7124
0    4089    7    6    2    4004    4020
0    4250    5    1    1    4247
0    4254    5    1    1    4251
0    4258    5    1    1    4255
0    4262    5    1    1    4259
0    4272    7    1    3    4189    4180    4247
0    4275    7    1    3    4193    4184    4251
0    4278    7    1    3    4212    4203    4255
0    4281    7    1    3    4216    4207    4259
0    4285    4    1    2    4283    4284
0    4288    4    1    2    4286    4287
0    4360    5    1    1    4356
0    4380    6    1    2    4369    89
0    4386    7    3    2    4356    4369
0    7442    5    1    1    7438
0    4609    5    1    1    4606
0    4613    5    1    1    4610
0    4617    5    1    1    4614
0    4621    5    1    1    4618
0    4624    4    1    2    4622    4623
0    4627    4    1    2    4625    4626
0    4629    7    1    3    4563    4554    4606
0    4632    7    1    3    4567    4558    4610
0    4635    7    1    3    4586    4577    4614
0    4638    7    1    3    4590    4581    4618
2    4836    1    2472
0    4949    6    2    2    4947    4948
0    4990    6    2    2    4988    4989
0    5020    6    1    2    5011    5018
0    5108    6    1    2    5099    5106
0    5590    6    1    2    5581    5588
0    5678    6    1    2    5669    5676
0    6084    5    1    1    6080
0    6094    5    1    1    6090
0    6104    5    1    1    6100
0    6142    5    1    1    6138
0    6152    5    1    1    6148
0    6162    5    1    1    6158
2    6206    1    2742
0    6220    5    1    1    6216
0    6230    5    1    1    6226
0    6240    5    1    1    6236
0    6328    5    1    1    6324
2    6294    1    2742
0    6308    5    1    1    6304
0    6318    5    1    1    6314
0    6362    6    2    2    6360    6361
0    6840    6    2    2    6817    6818
0    6848    6    2    2    6827    6828
0    6952    5    1    1    6948
0    6962    5    1    1    6958
0    6972    5    1    1    6968
0    7010    5    1    1    7006
0    7020    5    1    1    7016
0    7030    5    1    1    7026
0    7078    5    1    1    7074
0    7088    5    1    1    7084
0    7098    5    1    1    7094
0    7108    5    1    1    7104
0    7196    5    1    1    7192
0    7166    5    1    1    7162
0    7176    5    1    1    7172
0    7186    5    1    1    7182
0    7448    6    2    2    7446    7447
0    7458    6    2    2    7456    7457
0    254    7    1    2    3046    3249
0    260    7    1    2    3046    3249
0    1987    6    1    2    1985    1986
0    1994    6    1    2    1992    1993
0    2002    5    1    1    2001
0    962    7    2    2    933    924
0    1751    7    2    2    1730    1721
0    1990    6    1    2    1988    1989
0    1997    6    1    2    1995    1996
0    2499    5    1    1    2495
0    2536    7    1    2    2515    2487
0    5943    5    1    1    5937
0    2542    6    1    2    5937    5944
0    5951    5    1    1    5945
0    2545    6    1    2    5945    5952
0    5959    5    1    1    5953
0    2549    6    1    2    5953    5960
0    5967    5    1    1    5961
0    2552    6    1    2    5961    5968
0    2556    6    1    2    5969    5976
0    2560    6    1    2    5977    5984
0    2761    5    1    1    2757
0    2784    5    3    1    2780
0    2853    7    1    2    2749    2780
0    3135    5    1    1    3131
0    3146    5    1    1    3143
0    3163    7    1    2    3123    3143
0    3467    7    1    2    3453    3431
0    6645    5    1    1    6639
0    3470    6    1    2    6639    6646
0    6653    5    1    1    6647
0    3473    6    1    2    6647    6654
0    6661    5    1    1    6655
0    3477    6    1    2    6655    6662
0    6669    5    1    1    6663
0    3480    6    1    2    6663    6670
0    3484    6    1    2    6671    6678
0    3488    6    1    2    6679    6686
0    3601    7    1    3    3531    3536    3582
0    3604    7    1    3    3527    3540    3586
0    3607    7    1    3    3554    3559    3590
0    3610    7    1    3    3550    3563    3594
0    4032    5    2    1    4028
0    4090    7    1    2    4004    4028
0    4271    7    1    3    4184    4189    4250
0    4274    7    1    3    4180    4193    4254
0    4277    7    1    3    4207    4212    4258
0    4280    7    1    3    4203    4216    4262
0    4368    5    1    1    4364
0    4379    5    1    1    4376
0    4387    7    1    2    4356    4376
0    4628    7    1    3    4558    4563    4609
0    4631    7    1    3    4554    4567    4613
0    4634    7    1    3    4581    4586    4617
0    4637    7    1    3    4577    4590    4621
0    4841    3    2    5    2431    2518    2519    2520    2522
0    4849    3    2    4    2448    2523    2524    2526
0    4857    3    2    3    2465    2527    2529
0    4865    3    2    2    2481    2531
0    5021    6    2    2    5019    5020
0    5028    5    1    1    5024
0    5109    6    2    2    5107    5108
0    5116    5    1    1    5112
0    5369    6    2    2    1313    1310
0    5377    6    2    2    1319    1316
0    5385    6    2    2    1325    1322
0    5472    5    1    1    5468
0    5473    6    1    2    5468    5471
0    5530    5    1    1    5526
0    5531    6    1    2    5526    5529
0    5591    6    2    2    5589    5590
0    5598    5    1    1    5594
0    5679    6    2    2    5677    5678
0    5686    5    1    1    5682
0    6060    3    2    2    2768    2804
0    6074    5    1    1    6070
0    6118    5    2    1    2768
0    6132    5    1    1    6128
0    6176    3    2    4    2693    2795    2796    2797
0    6186    3    2    2    2801    2807
0    6196    3    2    5    2670    2788    2789    2790    2791
0    6268    5    1    1    6264
0    6269    6    1    2    6264    6267
0    6274    5    2    1    2801
0    6288    5    1    1    6284
0    6337    6    2    2    4288    4285
0    6829    6    2    2    3600    3597
0    6928    3    2    2    4017    4051
0    6942    5    1    1    6938
0    6986    5    2    1    4017
0    7000    5    1    1    6996
0    7048    5    1    1    7044
0    7049    6    1    2    7044    7047
0    7054    3    2    2    4048    4052
0    7068    5    1    1    7064
0    7136    5    1    1    7132
0    7137    6    1    2    7132    7135
0    7142    5    2    1    4048
0    7156    5    1    1    7152
0    7433    6    2    2    4627    4624
0    242    7    1    2    1982    1146
0    3151    6    1    2    3135    3127
0    257    7    1    5    89    4386    3156    3035    3249
0    263    7    1    5    89    4386    3156    3035    3249
0    266    7    1    2    1790    997
0    1991    5    1    1    1990
0    1998    5    1    1    1997
0    3489    6    1    2    3487    3488
0    371    6    1    2    4836    4839
0    4840    5    1    1    4836
0    2561    6    1    2    2559    2560
0    2532    7    3    2    2487    2508
0    2537    3    3    2    2495    2536
0    2541    6    1    2    5940    5943
0    2544    6    1    2    5948    5951
0    2548    6    1    2    5956    5959
0    2551    6    1    2    5964    5967
0    2557    6    1    2    2555    2556
0    2563    7    1    2    2508    4526
0    2577    6    1    2    2499    2491
0    2775    5    1    1    2771
0    2806    6    1    2    2771    4526
0    2808    6    1    2    2761    2753
0    2852    7    3    2    2749    2771
0    2854    3    3    2    2757    2853
0    6366    5    1    1    6362
0    4381    6    1    2    4368    4360
0    3164    3    3    2    3131    3163
0    3241    7    1    4    89    4386    3156    3035
0    3468    3    3    2    3437    3467
0    3469    6    1    2    6642    6645
0    3472    6    1    2    6650    6653
0    3476    6    1    2    6658    6661
0    3479    6    1    2    6666    6669
0    3485    6    1    2    3483    3484
0    3603    4    1    2    3601    3602
0    3606    4    1    2    3604    3605
0    3609    4    1    2    3607    3608
0    3612    4    1    2    3610    3611
0    6844    5    1    1    6840
0    6852    5    1    1    6848
0    4091    3    3    2    4010    4090
0    4273    4    1    2    4271    4272
0    4276    4    1    2    4274    4275
0    4279    4    1    2    4277    4278
0    4282    4    1    2    4280    4281
0    4382    7    2    2    4379    4380
0    4388    3    3    2    4364    4387
0    7452    5    1    1    7448
0    7462    5    1    1    7458
0    4630    4    1    2    4628    4629
0    4633    4    1    2    4631    4632
0    4636    4    1    2    4634    4635
0    4639    4    1    2    4637    4638
0    4955    5    1    1    4949
0    4958    6    1    2    4949    4956
0    4996    5    1    1    4990
0    4999    6    1    2    4990    4997
0    5474    6    1    2    5465    5472
0    5532    6    1    2    5523    5530
0    6210    5    1    1    6206
0    6270    6    1    2    6261    6268
0    6298    5    1    1    6294
0    7050    6    1    2    7041    7048
0    7138    6    1    2    7129    7136
0    3471    6    1    2    3469    3470
0    3478    6    1    2    3476    3477
0    3486    5    1    1    3485
0    372    6    1    2    4833    4840
0    2543    6    1    2    2541    2542
0    2550    6    1    2    2548    2549
0    2558    5    1    1    2557
0    4847    5    1    1    4841
0    387    6    1    2    4841    4848
0    4855    5    1    1    4849
0    390    6    1    2    4849    4856
0    4863    5    1    1    4857
0    393    6    1    2    4857    4864
0    4871    5    1    1    4865
0    396    6    1    2    4865    4872
0    965    5    1    1    962
0    5375    5    1    1    5369
0    1327    6    1    2    5369    5376
0    5383    5    1    1    5377
0    1330    6    1    2    5377    5384
0    5391    5    1    1    5385
0    1333    6    1    2    5385    5392
0    1754    5    1    1    1751
0    2546    6    1    2    2544    2545
0    2553    6    1    2    2551    2552
0    2564    3    6    2    2515    2563
0    2809    7    2    2    2784    2806
0    2813    7    2    2    2784    2775
0    6345    5    1    1    6337
0    2860    6    1    2    6337    6346
0    3474    6    1    2    3472    3473
0    3481    6    1    2    3479    3480
0    6835    5    1    1    6829
0    3614    6    1    2    6829    6836
0    4053    7    2    2    4032    4023
0    7441    5    1    1    7433
0    4516    6    1    2    7433    7442
0    4957    6    1    2    4952    4955
0    4998    6    1    2    4993    4996
0    5027    5    1    1    5021
0    5030    6    1    2    5021    5028
0    5115    5    1    1    5109
0    5118    6    1    2    5109    5116
0    5475    6    2    2    5473    5474
0    5533    6    2    2    5531    5532
0    5597    5    1    1    5591
0    5600    6    1    2    5591    5598
0    5685    5    1    1    5679
0    5688    6    1    2    5679    5686
0    6064    5    1    1    6060
0    6065    6    1    2    6060    6063
0    6122    5    1    1    6118
0    6123    6    1    2    6118    6121
0    6180    5    1    1    6176
0    6181    6    1    2    6176    6179
0    6190    5    1    1    6186
0    6200    5    1    1    6196
0    6271    6    2    2    6269    6270
0    6278    5    1    1    6274
0    6347    6    2    2    4276    4273
0    6357    6    2    2    4282    4279
0    6837    6    2    2    3606    3603
0    6845    6    2    2    3612    3609
0    6932    5    1    1    6928
0    6933    6    1    2    6928    6931
0    6990    5    1    1    6986
0    6991    6    1    2    6986    6989
0    7051    6    2    2    7049    7050
0    7058    5    1    1    7054
0    7139    6    2    2    7137    7138
0    7146    5    1    1    7142
0    7443    6    2    2    4639    4636
0    7453    6    2    2    4633    4630
0    243    7    1    3    3468    1974    1146
0    244    7    1    4    2537    3466    1974    1146
0    245    7    1    5    4526    2532    3466    1974    1146
0    255    7    1    3    3164    3035    3249
0    256    7    1    4    4388    3156    3035    3249
0    261    7    1    3    3164    3035    3249
0    262    7    1    4    4388    3156    3035    3249
0    267    7    1    3    4091    1788    997
0    268    7    1    4    2854    4089    1788    997
0    269    7    1    5    4526    2852    4089    1788    997
0    3475    5    1    1    3474
0    3482    5    1    1    3481
3    373    6    0    2    371    372
0    2547    5    1    1    2546
0    2554    5    1    1    2553
0    386    6    1    2    4844    4847
0    389    6    1    2    4852    4855
0    392    6    1    2    4860    4863
0    395    6    1    2    4868    4871
0    1326    6    1    2    5372    5375
0    1329    6    1    2    5380    5383
0    1332    6    1    2    5388    5391
0    1436    7    1    2    4091    1788
0    1440    7    1    3    2854    4089    1788
0    1445    7    1    4    4526    2852    4089    1788
0    1450    7    1    2    2854    4089
0    1454    7    1    3    4526    2852    4089
0    2859    6    1    2    6342    6345
0    4385    5    1    1    4382
0    3148    7    1    2    4382    4364
0    3239    7    1    2    3164    3035
0    3240    7    1    3    4388    3156    3035
0    3265    7    1    2    3468    1974
0    3267    7    1    3    2537    3466    1974
0    3270    7    1    4    4526    2532    3466    1974
0    3274    7    1    2    2537    3466
0    3277    7    1    3    4526    2532    3466
0    3613    6    1    2    6832    6835
0    4515    6    1    2    7438    7441
0    4959    6    2    2    4957    4958
0    5000    6    2    2    4998    4999
0    5029    6    1    2    5024    5027
0    5117    6    1    2    5112    5115
0    5599    6    1    2    5594    5597
0    5687    6    1    2    5682    5685
0    6066    6    1    2    6057    6064
0    6124    6    1    2    6115    6122
0    6182    6    1    2    6173    6180
0    6934    6    1    2    6925    6932
0    6992    6    1    2    6983    6990
3    246    3    0    5    241    242    243    244    245
3    258    3    0    5    3259    254    255    256    257
3    264    3    0    5    3259    260    261    262    263
3    270    3    0    5    265    266    267    268    269
0    375    7    1    2    2564    2543
0    378    7    1    2    2564    2550
0    381    7    1    2    2564    2558
0    384    7    1    2    2564    2406
3    388    6    0    2    386    387
3    391    6    0    2    389    390
3    394    6    0    2    392    393
3    397    6    0    2    395    396
0    1328    6    1    2    1326    1327
0    1331    6    1    2    1329    1330
0    1334    6    1    2    1332    1333
0    1447    3    2    4    1790    1436    1440    1445
0    1766    3    4    3    4091    1450    1454
0    2571    5    5    1    2564
0    2579    7    1    2    2577    2564
0    2812    5    1    1    2809
0    2816    5    1    1    2813
0    2851    7    1    2    2809    2757
0    2861    6    1    2    2859    2860
0    6355    5    1    1    6347
0    2863    6    1    2    6347    6356
0    6365    5    1    1    6357
0    2866    6    1    2    6357    6366
0    3147    7    1    2    4381    4385
0    3242    3    1    4    3046    3239    3240    3241
0    3271    3    6    4    1982    3265    3267    3270
0    3279    3    6    3    3468    3274    3277
0    3615    6    1    2    3613    3614
0    6843    5    1    1    6837
0    3617    6    1    2    6837    6844
0    6851    5    1    1    6845
0    3620    6    1    2    6845    6852
0    4056    5    1    1    4053
0    4517    6    1    2    4515    4516
0    7451    5    1    1    7443
0    4519    6    1    2    7443    7452
0    7461    5    1    1    7453
0    4522    6    1    2    7453    7462
0    5031    6    2    2    5029    5030
0    5119    6    2    2    5117    5118
0    5481    5    1    1    5475
0    5484    6    1    2    5475    5482
0    5539    5    1    1    5533
0    5542    6    1    2    5533    5540
0    5601    6    2    2    5599    5600
0    5689    6    2    2    5687    5688
0    6067    6    2    2    6065    6066
0    6125    6    2    2    6123    6124
0    6183    6    2    2    6181    6182
0    6277    5    1    1    6271
0    6280    6    1    2    6271    6278
0    6935    6    2    2    6933    6934
0    6993    6    2    2    6991    6992
0    7057    5    1    1    7051
0    7060    6    1    2    7051    7058
0    7145    5    1    1    7139
0    7148    6    1    2    7139    7146
0    4968    6    1    2    4959    4966
0    5009    6    1    2    5000    5007
0    2850    7    1    2    2808    2812
0    2862    6    1    2    6352    6355
0    2865    6    1    2    6362    6365
0    3149    3    1    2    3147    3148
0    3243    6    1    2    3228    3242
0    3616    6    1    2    6840    6843
0    3619    6    1    2    6848    6851
0    4518    6    1    2    7448    7451
0    4521    6    1    2    7458    7461
0    4965    5    1    1    4959
0    5006    5    1    1    5000
0    5483    6    1    2    5478    5481
0    5541    6    1    2    5536    5539
0    6279    6    1    2    6274    6277
0    7059    6    1    2    7054    7057
0    7147    6    1    2    7142    7145
0    374    7    1    2    2547    2571
0    377    7    1    2    2554    2571
0    380    7    1    2    2561    2571
0    383    7    1    2    2400    2571
0    955    6    1    2    920    1447
0    4967    6    1    2    4962    4965
0    5008    6    1    2    5003    5006
2    975    1    1447
0    1136    7    1    5    3271    1093    1055    1074    1038
0    1140    7    1    4    3271    1093    1055    1074
0    1143    7    1    3    3271    1093    1074
0    1145    7    1    2    3271    1093
0    1160    7    1    2    1122    3271
0    1771    5    3    1    1766
0    1964    7    1    5    3279    1921    1885    1903    1869
0    1968    7    1    4    3279    1921    1885    1903
0    1971    7    1    3    3279    1921    1903
0    1973    7    1    2    3279    1921
0    2007    7    1    2    1950    3279
0    2578    7    1    2    2495    2571
0    2864    6    1    2    2862    2863
0    2867    6    1    2    2865    2866
0    3150    6    1    2    3136    3149
0    3245    7    2    2    3238    3243
0    3618    6    1    2    3616    3617
0    3621    6    1    2    3619    3620
0    4067    3    4    2    2850    2851
0    4520    6    1    2    4518    4519
0    4523    6    1    2    4521    4522
2    4713    1    3279
2    4753    1    3271
0    5037    5    1    1    5031
0    5040    6    1    2    5031    5038
0    5125    5    1    1    5119
0    5128    6    1    2    5119    5126
0    5485    6    2    2    5483    5484
0    5543    6    2    2    5541    5542
0    5607    5    1    1    5601
0    5610    6    1    2    5601    5608
0    5695    5    1    1    5689
0    5698    6    1    2    5689    5696
0    6073    5    1    1    6067
0    6076    6    1    2    6067    6074
0    6131    5    1    1    6125
0    6134    6    1    2    6125    6132
0    6189    5    1    1    6183
0    6192    6    1    2    6183    6190
0    6281    6    2    2    6279    6280
0    6941    5    1    1    6935
0    6944    6    1    2    6935    6942
0    6999    5    1    1    6993
0    7002    6    1    2    6993    7000
0    7061    6    2    2    7059    7060
0    7149    6    2    2    7147    7148
3    376    3    0    2    374    375
3    379    3    0    2    377    378
3    382    3    0    2    380    381
3    385    3    0    2    383    384
0    958    7    2    2    933    955
0    967    6    2    2    4967    4968
0    971    6    2    2    5008    5009
0    1161    3    4    2    1129    1160
0    2008    3    5    2    1957    2007
0    2580    3    6    2    2578    2579
0    2868    7    2    4    1331    2861    2864    2867
0    3152    7    2    2    3146    3150
0    4443    7    2    4    1328    1334    3618    3621
0    4524    7    2    4    3615    4517    4520    4523
0    4721    3    2    5    1880    1960    1961    1962    1964
0    4729    3    2    4    1897    1965    1966    1968
0    4737    3    2    3    1914    1969    1971
0    4745    3    2    2    1929    1973
0    4761    3    2    5    1050    1132    1133    1134    1136
0    4769    3    2    4    1068    1137    1138    1140
0    4777    3    2    3    1086    1141    1143
0    4785    3    2    2    1102    1145
0    5039    6    1    2    5034    5037
0    5127    6    1    2    5122    5125
0    5609    6    1    2    5604    5607
0    5697    6    1    2    5692    5695
0    6075    6    1    2    6070    6073
0    6133    6    1    2    6128    6131
0    6191    6    1    2    6186    6189
0    6943    6    1    2    6938    6941
0    7001    6    1    2    6996    6999
0    3248    5    1    1    3245
0    248    7    1    2    3245    3223
0    4719    5    1    1    4713
0    294    6    1    2    4713    4720
0    4759    5    1    1    4753
0    323    6    1    2    4753    4760
0    980    5    3    1    975
0    4072    5    3    1    4067
0    5041    6    2    2    5039    5040
0    5129    6    2    2    5127    5128
0    5491    5    1    1    5485
0    5494    6    1    2    5485    5492
0    5549    5    1    1    5543
0    5552    6    1    2    5543    5550
0    5611    6    2    2    5609    5610
0    5699    6    2    2    5697    5698
0    6077    6    2    2    6075    6076
0    6135    6    2    2    6133    6134
0    6193    6    2    2    6191    6192
0    6287    5    1    1    6281
0    6290    6    1    2    6281    6288
0    6945    6    2    2    6943    6944
0    7003    6    2    2    7001    7002
0    7067    5    1    1    7061
0    7070    6    1    2    7061    7068
0    7155    5    1    1    7149
0    7158    6    1    2    7149    7156
0    247    7    1    2    3244    3248
0    3155    5    1    1    3152
0    251    7    1    2    3152    3131
0    272    7    1    2    1176    1161
0    961    5    1    1    958
0    275    7    1    2    958    908
0    293    6    1    2    4716    4719
0    297    7    1    2    2008    1987
0    300    7    1    2    2008    1994
0    303    7    1    2    2008    2002
0    306    7    1    2    2008    1856
0    4727    5    1    1    4721
0    309    6    1    2    4721    4728
0    4735    5    1    1    4729
0    312    6    1    2    4729    4736
0    4743    5    1    1    4737
0    315    6    1    2    4737    4744
0    4751    5    1    1    4745
0    318    6    1    2    4745    4752
0    322    6    1    2    4756    4759
0    4767    5    1    1    4761
0    326    6    1    2    4761    4768
0    4775    5    1    1    4769
0    329    6    1    2    4769    4776
0    4783    5    1    1    4777
0    332    6    1    2    4777    4784
0    4791    5    1    1    4785
0    335    6    1    2    4785    4792
3    412    5    0    1    4443
3    414    5    0    1    4524
3    416    5    0    1    2868
0    2881    7    1    3    4443    4524    2868
0    993    7    1    3    971    962    975
0    994    7    1    3    967    965    975
0    1166    5    3    1    1161
0    1171    7    1    2    1161    1155
0    1174    7    1    2    1161    1023
0    2014    5    4    1    2008
0    3459    7    1    5    2580    3417    3381    3399    3365
0    3462    7    1    4    2580    3417    3381    3399
0    3464    7    1    3    2580    3417    3399
0    3465    7    1    2    2580    3417
0    3490    7    1    2    3446    2580
2    4793    1    2580
0    5493    6    1    2    5488    5491
0    5551    6    1    2    5546    5549
0    6289    6    1    2    6284    6287
0    7069    6    1    2    7064    7067
0    7157    6    1    2    7152    7155
3    249    3    0    2    247    248
0    250    7    1    2    3151    3155
0    274    7    1    2    957    961
3    295    6    0    2    293    294
0    308    6    1    2    4724    4727
0    311    6    1    2    4732    4735
0    314    6    1    2    4740    4743
0    317    6    1    2    4748    4751
3    324    6    0    2    322    323
0    325    6    1    2    4764    4767
0    328    6    1    2    4772    4775
0    331    6    1    2    4780    4783
0    334    6    1    2    4788    4791
0    417    7    1    3    2876    2878    2881
0    991    7    1    3    971    933    980
0    992    7    1    3    967    929    980
0    3491    3    5    2    3453    3490
0    4801    3    2    5    3376    3456    3457    3458    3459
0    4809    3    2    4    3393    3460    3461    3462
0    4817    3    2    3    3410    3463    3464
0    4825    3    2    2    3425    3465
0    5047    5    1    1    5041
0    5050    6    1    2    5041    5048
0    5135    5    1    1    5129
0    5138    6    1    2    5129    5136
0    5495    6    2    2    5493    5494
0    5553    6    2    2    5551    5552
0    5617    5    1    1    5611
0    5620    6    1    2    5611    5618
0    5705    5    1    1    5699
0    5708    6    1    2    5699    5706
0    6083    5    1    1    6077
0    6086    6    1    2    6077    6084
0    6141    5    1    1    6135
0    6144    6    1    2    6135    6142
0    6199    5    1    1    6193
0    6202    6    1    2    6193    6200
0    6291    6    2    2    6289    6290
0    6951    5    1    1    6945
0    6954    6    1    2    6945    6952
0    7009    5    1    1    7003
0    7012    6    1    2    7003    7010
0    7071    6    2    2    7069    7070
0    7159    6    2    2    7157    7158
3    252    3    0    2    250    251
0    271    7    1    2    1117    1166
3    276    3    0    2    274    275
0    296    7    1    2    1991    2014
0    299    7    1    2    1998    2014
0    302    7    1    2    2005    2014
0    305    7    1    2    1850    2014
3    310    6    0    2    308    309
3    313    6    0    2    311    312
3    316    6    0    2    314    315
3    319    6    0    2    317    318
3    327    6    0    2    325    326
3    330    6    0    2    328    329
3    333    6    0    2    331    332
3    336    6    0    2    334    335
0    4799    5    1    1    4793
0    343    6    1    2    4793    4800
3    418    5    0    1    417
0    1170    7    1    2    1158    1166
0    1173    7    1    2    1019    1166
0    5049    6    1    2    5044    5047
0    5137    6    1    2    5132    5135
0    5167    3    2    4    991    992    993    994
0    5619    6    1    2    5614    5617
0    5707    6    1    2    5702    5705
0    6085    6    1    2    6080    6083
0    6143    6    1    2    6138    6141
0    6201    6    1    2    6196    6199
0    6953    6    1    2    6948    6951
0    7011    6    1    2    7006    7009
3    273    3    0    2    271    272
3    298    3    0    2    296    297
3    301    3    0    2    299    300
3    304    3    0    2    302    303
3    307    3    0    2    305    306
0    342    6    1    2    4796    4799
0    346    7    1    2    3491    3471
0    349    7    1    2    3491    3478
0    352    7    1    2    3491    3486
0    355    7    1    2    3491    3350
0    4807    5    1    1    4801
0    358    6    1    2    4801    4808
0    4815    5    1    1    4809
0    361    6    1    2    4809    4816
0    4823    5    1    1    4817
0    364    6    1    2    4817    4824
0    4831    5    1    1    4825
0    367    6    1    2    4825    4832
0    1172    3    2    2    1170    1171
0    1175    3    2    2    1173    1174
0    3497    5    4    1    3491
0    5051    6    2    2    5049    5050
0    5139    6    2    2    5137    5138
0    5501    5    1    1    5495
0    5504    6    1    2    5495    5502
0    5559    5    1    1    5553
0    5562    6    1    2    5553    5560
0    5621    6    2    2    5619    5620
0    5709    6    2    2    5707    5708
0    6087    6    2    2    6085    6086
0    6145    6    2    2    6143    6144
0    6203    6    2    2    6201    6202
0    6297    5    1    1    6291
0    6300    6    1    2    6291    6298
0    6955    6    2    2    6953    6954
0    7013    6    2    2    7011    7012
0    7077    5    1    1    7071
0    7080    6    1    2    7071    7078
0    7165    5    1    1    7159
0    7168    6    1    2    7159    7166
3    344    6    0    2    342    343
0    357    6    1    2    4804    4807
0    360    6    1    2    4812    4815
0    363    6    1    2    4820    4823
0    366    6    1    2    4828    4831
0    5173    5    1    1    5167
3    422    1    0    1    1172
3    469    1    0    1    1172
3    419    1    0    1    1175
3    471    1    0    1    1175
0    5503    6    1    2    5498    5501
0    5561    6    1    2    5556    5559
0    6299    6    1    2    6294    6297
0    7079    6    1    2    7074    7077
0    7167    6    1    2    7162    7165
0    345    7    1    2    3475    3497
0    348    7    1    2    3482    3497
0    351    7    1    2    3489    3497
0    354    7    1    2    3344    3497
3    359    6    0    2    357    358
3    362    6    0    2    360    361
3    365    6    0    2    363    364
3    368    6    0    2    366    367
0    5057    5    1    1    5051
0    5060    6    1    2    5051    5058
0    5145    5    1    1    5139
0    5148    6    1    2    5139    5146
0    5505    6    2    2    5503    5504
0    5563    6    2    2    5561    5562
0    5627    5    1    1    5621
0    5630    6    1    2    5621    5628
0    5715    5    1    1    5709
0    5718    6    1    2    5709    5716
0    6093    5    1    1    6087
0    6096    6    1    2    6087    6094
0    6151    5    1    1    6145
0    6154    6    1    2    6145    6152
0    6209    5    1    1    6203
0    6212    6    1    2    6203    6210
0    6301    6    2    2    6299    6300
0    6961    5    1    1    6955
0    6964    6    1    2    6955    6962
0    7019    5    1    1    7013
0    7022    6    1    2    7013    7020
0    7081    6    2    2    7079    7080
0    7169    6    2    2    7167    7168
3    347    3    0    2    345    346
3    350    3    0    2    348    349
3    353    3    0    2    351    352
3    356    3    0    2    354    355
0    5059    6    1    2    5054    5057
0    5147    6    1    2    5142    5145
0    5629    6    1    2    5624    5627
0    5717    6    1    2    5712    5715
0    6095    6    1    2    6090    6093
0    6153    6    1    2    6148    6151
0    6211    6    1    2    6206    6209
0    6963    6    1    2    6958    6961
0    7021    6    1    2    7016    7019
0    5061    6    2    2    5059    5060
0    5149    6    2    2    5147    5148
0    5511    5    1    1    5505
0    5514    6    1    2    5505    5512
0    5569    5    1    1    5563
0    5572    6    1    2    5563    5570
0    5631    6    2    2    5629    5630
0    5719    6    2    2    5717    5718
0    6097    6    2    2    6095    6096
0    6155    6    2    2    6153    6154
0    6213    6    2    2    6211    6212
0    6307    5    1    1    6301
0    6310    6    1    2    6301    6308
0    6965    6    2    2    6963    6964
0    7023    6    2    2    7021    7022
0    7087    5    1    1    7081
0    7090    6    1    2    7081    7088
0    7175    5    1    1    7169
0    7178    6    1    2    7169    7176
0    5513    6    1    2    5508    5511
0    5571    6    1    2    5566    5569
0    6309    6    1    2    6304    6307
0    7089    6    1    2    7084    7087
0    7177    6    1    2    7172    7175
0    5067    5    1    1    5061
0    5070    6    1    2    5061    5068
0    5155    5    1    1    5149
0    5158    6    1    2    5149    5156
0    5515    6    2    2    5513    5514
0    5573    6    2    2    5571    5572
0    5637    5    1    1    5631
0    5640    6    1    2    5631    5638
0    5725    5    1    1    5719
0    5728    6    1    2    5719    5726
0    6103    5    1    1    6097
0    6106    6    1    2    6097    6104
0    6161    5    1    1    6155
0    6164    6    1    2    6155    6162
0    6219    5    1    1    6213
0    6222    6    1    2    6213    6220
0    6311    6    2    2    6309    6310
0    6971    5    1    1    6965
0    6974    6    1    2    6965    6972
0    7029    5    1    1    7023
0    7032    6    1    2    7023    7030
0    7091    6    2    2    7089    7090
0    7179    6    2    2    7177    7178
0    5069    6    1    2    5064    5067
0    5157    6    1    2    5152    5155
0    5639    6    1    2    5634    5637
0    5727    6    1    2    5722    5725
0    6105    6    1    2    6100    6103
0    6163    6    1    2    6158    6161
0    6221    6    1    2    6216    6219
0    6973    6    1    2    6968    6971
0    7031    6    1    2    7026    7029
0    5521    5    1    1    5515
0    1756    6    1    2    5515    5522
0    5579    5    1    1    5573
0    1761    6    1    2    5573    5580
0    5071    6    2    2    5069    5070
0    5159    6    2    2    5157    5158
0    5641    6    2    2    5639    5640
0    5729    6    2    2    5727    5728
0    6107    6    2    2    6105    6106
0    6165    6    2    2    6163    6164
0    6223    6    2    2    6221    6222
0    6317    5    1    1    6311
0    6320    6    1    2    6311    6318
0    6975    6    2    2    6973    6974
0    7033    6    2    2    7031    7032
0    7097    5    1    1    7091
0    7100    6    1    2    7091    7098
0    7185    5    1    1    7179
0    7188    6    1    2    7179    7186
0    1755    6    1    2    5518    5521
0    1760    6    1    2    5576    5579
0    6319    6    1    2    6314    6317
0    7099    6    1    2    7094    7097
0    7187    6    1    2    7182    7185
0    1757    6    2    2    1755    1756
0    1762    6    2    2    1760    1761
0    6113    5    1    1    6107
0    2818    6    1    2    6107    6114
0    6171    5    1    1    6165
0    2823    6    1    2    6165    6172
0    6981    5    1    1    6975
0    4058    6    1    2    6975    6982
0    7039    5    1    1    7033
0    4063    6    1    2    7033    7040
0    5077    5    1    1    5071
0    5080    6    1    2    5071    5078
0    5165    5    1    1    5159
0    5090    6    1    2    5159    5166
0    5647    5    1    1    5641
0    5650    6    1    2    5641    5648
0    5735    5    1    1    5729
0    5660    6    1    2    5729    5736
0    6229    5    1    1    6223
0    6232    6    1    2    6223    6230
0    6321    6    2    2    6319    6320
0    7101    6    2    2    7099    7100
0    7189    6    2    2    7187    7188
0    2817    6    1    2    6110    6113
0    2822    6    1    2    6168    6171
0    4057    6    1    2    6978    6981
0    4062    6    1    2    7036    7039
0    5079    6    1    2    5074    5077
0    5089    6    1    2    5162    5165
0    5649    6    1    2    5644    5647
0    5659    6    1    2    5732    5735
0    6231    6    1    2    6226    6229
0    1782    7    1    3    1762    1730    1771
0    1783    7    1    3    1757    1726    1771
0    1784    7    1    3    1762    1751    1766
0    1785    7    1    3    1757    1754    1766
0    2819    6    2    2    2817    2818
0    2824    6    2    2    2822    2823
0    4059    6    2    2    4057    4058
0    4064    6    2    2    4062    4063
0    5081    6    2    2    5079    5080
0    5091    6    2    2    5089    5090
0    5651    6    2    2    5649    5650
0    5661    6    2    2    5659    5660
0    6233    6    2    2    6231    6232
0    6327    5    1    1    6321
0    6252    6    1    2    6321    6328
0    7107    5    1    1    7101
0    7110    6    1    2    7101    7108
0    7195    5    1    1    7189
0    7120    6    1    2    7189    7196
0    5737    3    2    4    1782    1783    1784    1785
0    6251    6    1    2    6324    6327
0    7109    6    1    2    7104    7107
0    7119    6    1    2    7192    7195
0    5087    5    1    1    5081
0    985    6    1    2    5081    5088
0    5097    5    1    1    5091
0    988    6    1    2    5091    5098
0    5657    5    1    1    5651
0    1776    6    1    2    5651    5658
0    5667    5    1    1    5661
0    1779    6    1    2    5661    5668
0    2844    7    1    3    2824    2784    2833
0    2845    7    1    3    2819    2780    2833
0    2846    7    1    3    2824    2813    2828
0    2847    7    1    3    2819    2816    2828
0    4083    7    1    3    4064    4032    4072
0    4084    7    1    3    4059    4028    4072
0    4085    7    1    3    4064    4053    4067
0    4086    7    1    3    4059    4056    4067
0    6239    5    1    1    6233
0    6242    6    1    2    6233    6240
0    6253    6    2    2    6251    6252
0    7111    6    2    2    7109    7110
0    7121    6    2    2    7119    7120
0    984    6    1    2    5084    5087
0    987    6    1    2    5094    5097
0    1775    6    1    2    5654    5657
0    1778    6    1    2    5664    5667
0    5743    5    1    1    5737
0    6241    6    1    2    6236    6239
0    6329    3    2    4    2844    2845    2846    2847
0    7197    3    2    4    4083    4084    4085    4086
0    986    6    1    2    984    985
0    989    6    1    2    987    988
0    1777    6    1    2    1775    1776
0    1780    6    1    2    1778    1779
0    6259    5    1    1    6253
0    2841    6    1    2    6253    6260
0    7117    5    1    1    7111
0    4077    6    1    2    7111    7118
0    7127    5    1    1    7121
0    4080    6    1    2    7121    7128
0    6243    6    2    2    6241    6242
0    990    5    1    1    989
0    996    7    1    2    975    986
0    1781    5    1    1    1780
0    1787    7    1    2    1766    1777
0    2840    6    1    2    6256    6259
0    6335    5    1    1    6329
0    4076    6    1    2    7114    7117
0    4079    6    1    2    7124    7127
0    7203    5    1    1    7197
0    995    7    1    2    990    980
0    1786    7    1    2    1781    1771
0    6249    5    1    1    6243
0    2838    6    1    2    6243    6250
0    2842    6    1    2    2840    2841
0    4078    6    1    2    4076    4077
0    4081    6    1    2    4079    4080
0    2837    6    1    2    6246    6249
0    2843    5    1    1    2842
0    4082    5    1    1    4081
0    4088    7    1    2    4067    4078
0    5170    3    2    2    995    996
0    5740    3    2    2    1786    1787
0    2839    6    1    2    2837    2838
0    2848    7    1    2    2843    2833
0    4087    7    1    2    4082    4072
0    1791    6    1    2    5740    5743
0    1003    6    1    2    5170    5173
0    5174    5    1    1    5170
0    5744    5    1    1    5740
0    2849    7    1    2    2828    2839
0    7200    3    2    2    4087    4088
0    1792    6    1    2    5737    5744
0    1004    6    1    2    5167    5174
0    6332    3    2    2    2848    2849
0    320    6    1    2    1791    1792
0    337    6    1    2    1003    1004
0    4092    6    1    2    7200    7203
0    7204    5    1    1    7200
3    321    5    0    1    320
3    338    5    0    1    337
0    4093    6    1    2    7197    7204
0    2855    6    1    2    6332    6335
0    6336    5    1    1    6332
0    369    6    1    2    4092    4093
0    2856    6    1    2    6329    6336
3    370    5    0    1    369
0    398    6    1    2    2855    2856
3    399    5    0    1    398
3    339    0    0    0
